test of pipo adder and piso
.lib '/class/ece482/gpdk045_mos' SS

$The following parameter can be modified.
.param TCK = 0.430n

$The following parameters cannot be modified.
.param trf_ck = 5p
.param trf_ip_reset = 50p
.param CK_pw = 0.5*TCK
.param reset_delay = 0
.param reset_delay2 = 40*TCK
.param reset_pw = 0.9n
.param reset_pw2 = 5n
.param sim_end = 80*TCK
.param input_delay = 0.5n
.param input_pw = 4*TCK
.param input_delay_re = 10*TCK
.param input_delay_re2 = reset_pw2+4*TCK

$Clock Buffer - You will clk_out as your clock signal
mnm1 clk_out net10 vss vss g45n1svt L=45e-9 W=960e-9 AD=134.4e-15 AS=134.4e-15 PD=2.2e-6 PS=2.2e-6 NRD=145.833e-3 NRS=145.833e-3 M=1
mnm0 net10 CK vss vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm1 clk_out net10 vdd vdd g45p1svt L=45e-9 W=1.92e-6 AD=268.8e-15 AS=268.8e-15 PD=4.12e-6 PS=4.12e-6 NRD=72.9167e-3 NRS=72.9167e-3 M=1
mpm0 net10 CK vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1

vX3 x3 0 PWL(0 0 'input_delay+0*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+0*input_pw' 1.1 'input_delay+1*trf_ip_reset+1*input_pw' 1.1 'input_delay+2*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+2*input_pw' 0 'input_delay+3*trf_ip_reset+2*input_pw' 1.1 'input_delay+3*trf_ip_reset+3*input_pw' 1.1  'input_delay+4*trf_ip_reset+3*input_pw' 0 'input_delay+4*trf_ip_reset+4*input_pw' 0 'input_delay+5*trf_ip_reset+4*input_pw' 1.1 'input_delay+5*trf_ip_reset+5*input_pw' 1.1 'input_delay+6*trf_ip_reset+5*input_pw' 0 'input_delay+6*trf_ip_reset+6*input_pw' 0 'input_delay+7*trf_ip_reset+6*input_pw' 1.1 'input_delay+7*trf_ip_reset+7*input_pw' 1.1 'input_delay+8*trf_ip_reset+7*input_pw' 0 'input_delay+8*trf_ip_reset+8*input_pw' 0  'input_delay+8*trf_ip_reset+8*input_pw+input_delay_re' 0 'input_delay+9*trf_ip_reset+8*input_pw+input_delay_re' 1.1 'input_delay+9*trf_ip_reset+9*input_pw+input_delay_re' 1.1 'input_delay+10*trf_ip_reset+9*input_pw+input_delay_re' 0 'input_delay+10*trf_ip_reset+9*input_pw+input_delay_re++input_delay_re2' 0 'input_delay+11*trf_ip_reset+9*input_pw+input_delay_re++input_delay_re2' 1.1 'input_delay+11*trf_ip_reset+10*input_pw+input_delay_re++input_delay_re2' 1.1 'input_delay+12*trf_ip_reset+10*input_pw+input_delay_re++input_delay_re2' 0 sim_end 0)
vX2 x2 0 PWL(0 0 'input_delay+0*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+0*input_pw' 1.1 'input_delay+1*trf_ip_reset+1*input_pw' 1.1 'input_delay+2*trf_ip_reset+1*input_pw' 1.1 'input_delay+2*trf_ip_reset+2*input_pw' 1.1 'input_delay+3*trf_ip_reset+2*input_pw' 0 'input_delay+3*trf_ip_reset+3*input_pw' 0  'input_delay+4*trf_ip_reset+3*input_pw' 0 'input_delay+4*trf_ip_reset+4*input_pw' 0 'input_delay+5*trf_ip_reset+4*input_pw' 1.1 'input_delay+5*trf_ip_reset+5*input_pw' 1.1 'input_delay+6*trf_ip_reset+5*input_pw' 1.1 'input_delay+6*trf_ip_reset+6*input_pw' 1.1 'input_delay+7*trf_ip_reset+6*input_pw' 0 'input_delay+7*trf_ip_reset+7*input_pw' 0 'input_delay+8*trf_ip_reset+7*input_pw' 0 'input_delay+8*trf_ip_reset+8*input_pw' 0 sim_end 0)
vX1 x1 0 PWL(0 0 'input_delay+0*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+0*input_pw' 1.1 'input_delay+1*trf_ip_reset+1*input_pw' 1.1 'input_delay+2*trf_ip_reset+1*input_pw' 1.1 'input_delay+2*trf_ip_reset+2*input_pw' 1.1 'input_delay+3*trf_ip_reset+2*input_pw' 1.1 'input_delay+3*trf_ip_reset+3*input_pw' 1.1  'input_delay+4*trf_ip_reset+3*input_pw' 1.1 'input_delay+4*trf_ip_reset+4*input_pw' 1.1 'input_delay+5*trf_ip_reset+4*input_pw' 0 'input_delay+5*trf_ip_reset+5*input_pw' 0 'input_delay+6*trf_ip_reset+5*input_pw' 0 'input_delay+6*trf_ip_reset+6*input_pw' 0 'input_delay+7*trf_ip_reset+6*input_pw' 0 'input_delay+7*trf_ip_reset+7*input_pw' 0 'input_delay+8*trf_ip_reset+7*input_pw' 0 'input_delay+8*trf_ip_reset+8*input_pw' 0 sim_end 0)
vX0 x0 0 PWL(0 0 'input_delay+0*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+0*input_pw' 1.1 'input_delay+1*trf_ip_reset+1*input_pw' 1.1 'input_delay+2*trf_ip_reset+1*input_pw' 1.1 'input_delay+2*trf_ip_reset+2*input_pw' 1.1 'input_delay+3*trf_ip_reset+2*input_pw' 1.1 'input_delay+3*trf_ip_reset+3*input_pw' 1.1  'input_delay+4*trf_ip_reset+3*input_pw' 1.1 'input_delay+4*trf_ip_reset+4*input_pw' 1.1 'input_delay+5*trf_ip_reset+4*input_pw' 1.1 'input_delay+5*trf_ip_reset+5*input_pw' 1.1 'input_delay+6*trf_ip_reset+5*input_pw' 1.1 'input_delay+6*trf_ip_reset+6*input_pw' 1.1 'input_delay+7*trf_ip_reset+6*input_pw' 1.1 'input_delay+7*trf_ip_reset+7*input_pw' 1.1 'input_delay+8*trf_ip_reset+7*input_pw' 1.1 'input_delay+8*trf_ip_reset+8*input_pw' 1.1 sim_end 1.1)
vY3 y3 0 PWL(0 0 'input_delay+0*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+2*input_pw' 0 'input_delay+3*trf_ip_reset+2*input_pw' 0 'input_delay+3*trf_ip_reset+3*input_pw' 0  'input_delay+4*trf_ip_reset+3*input_pw' 0 'input_delay+4*trf_ip_reset+4*input_pw' 0 'input_delay+5*trf_ip_reset+4*input_pw' 1.1 'input_delay+5*trf_ip_reset+5*input_pw' 1.1 'input_delay+6*trf_ip_reset+5*input_pw' 1.1 'input_delay+6*trf_ip_reset+6*input_pw' 1.1 'input_delay+7*trf_ip_reset+6*input_pw' 1.1 'input_delay+7*trf_ip_reset+7*input_pw' 1.1 'input_delay+8*trf_ip_reset+7*input_pw' 1.1 'input_delay+8*trf_ip_reset+8*input_pw' 1.1 sim_end 1.1)
vY2 y2 0 PWL(0 0 'input_delay+0*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+2*input_pw' 0 'input_delay+3*trf_ip_reset+2*input_pw' 0 'input_delay+3*trf_ip_reset+3*input_pw' 0  'input_delay+4*trf_ip_reset+3*input_pw' 0 'input_delay+4*trf_ip_reset+4*input_pw' 0 'input_delay+5*trf_ip_reset+4*input_pw' 1.1 'input_delay+5*trf_ip_reset+5*input_pw' 1.1 'input_delay+6*trf_ip_reset+5*input_pw' 1.1 'input_delay+6*trf_ip_reset+6*input_pw' 1.1 'input_delay+7*trf_ip_reset+6*input_pw' 1.1 'input_delay+7*trf_ip_reset+7*input_pw' 1.1 'input_delay+8*trf_ip_reset+7*input_pw' 1.1 'input_delay+8*trf_ip_reset+8*input_pw' 1.1 sim_end 1.1)
vY1 y1 0 PWL(0 0 'input_delay+0*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+2*input_pw' 0 'input_delay+3*trf_ip_reset+2*input_pw' 0 'input_delay+3*trf_ip_reset+3*input_pw' 0  'input_delay+4*trf_ip_reset+3*input_pw' 0 'input_delay+4*trf_ip_reset+4*input_pw' 0 'input_delay+5*trf_ip_reset+4*input_pw' 1.1 'input_delay+5*trf_ip_reset+5*input_pw' 1.1 'input_delay+6*trf_ip_reset+5*input_pw' 1.1 'input_delay+6*trf_ip_reset+6*input_pw' 1.1 'input_delay+7*trf_ip_reset+6*input_pw' 1.1 'input_delay+7*trf_ip_reset+7*input_pw' 1.1 'input_delay+8*trf_ip_reset+7*input_pw' 1.1 'input_delay+8*trf_ip_reset+8*input_pw' 1.1 sim_end 1.1)
vY0 y0 0 PWL(0 0 'input_delay+0*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+2*input_pw' 0 'input_delay+3*trf_ip_reset+2*input_pw' 0 'input_delay+3*trf_ip_reset+3*input_pw' 0  'input_delay+4*trf_ip_reset+3*input_pw' 0 'input_delay+4*trf_ip_reset+4*input_pw' 0 'input_delay+5*trf_ip_reset+4*input_pw' 1.1 'input_delay+5*trf_ip_reset+5*input_pw' 1.1 'input_delay+6*trf_ip_reset+5*input_pw' 1.1 'input_delay+6*trf_ip_reset+6*input_pw' 1.1 'input_delay+7*trf_ip_reset+6*input_pw' 1.1 'input_delay+7*trf_ip_reset+7*input_pw' 1.1 'input_delay+8*trf_ip_reset+7*input_pw' 1.1 'input_delay+8*trf_ip_reset+8*input_pw' 1.1 sim_end 1.1)

vCK CK 0 pulse(0 1.1 trf_ck trf_ck trf_ck CK_pw TCK)
vReset reset 0 PWL(0 1.1 reset_delay 1.1 'reset_delay+trf_ip_reset' 1.1 'reset_delay+reset_pw+trf_ip_reset' 1.1 'reset_delay+reset_pw+2*trf_ip_reset' 0 'reset_delay+reset_pw+2*trf_ip_reset+reset_delay2' 0 'reset_delay+reset_pw+3*trf_ip_reset+reset_delay2' 1.1 'reset_delay+reset_pw+reset_pw2+3*trf_ip_reset+reset_delay2' 1.1 'reset_delay+reset_pw+reset_pw2+4*trf_ip_reset+reset_delay2' 0 sim_end 0)

vVDDIO VDDIO 0 1.8
vVDD VDD 0 1.1
vVSS VSS 0 0

.tran 0 sim_end

.option post
c1 vdd vss 1.73361e-15
c2 chipdriverout vss 654.947e-18
c3 piso_out vss 424.755e-18
c4 reset vss 80.1019e-18
c5 shift vss 139.638e-18
c6 vddio vss 315.356e-18
c7 x0 vss 23.2767e-18
c8 x1 vss 37.4114e-18
c9 y0 vss 20.1309e-18
c10 y1 vss 32.8957e-18
c11 y2 vss 27.4975e-18
c12 y3 vss 28.3605e-18
c13 clk_out vss 128.156e-18
c14 piso_outinv vss 29.5964e-18
c15 bufin vss 38.4996e-18
c16 i5__clk_buf vss 24.8505e-18
c17 i5__r2 vss 38.8531e-18
c18 i5__r1 vss 146.445e-18
c19 i5__r0 vss 47.4403e-18
c20 i5__clk4 vss 30.8437e-18
c21 i5__i8__net2 vss 22.1376e-18
c22 i5__i8__net1 vss 46.1767e-18
c23 i5__i8__net4 vss 28.7577e-18
c24 i5__i8__net5 vss 46.3619e-18
c25 i5__i8__i10__net22 vss 46.648e-18
c26 i5__i8__i10__net23 vss 113.303e-21
c27 i5__i8__i10__net24 vss 49.9317e-18
c28 i5__i8__i10__net21 vss 101.594e-21
c29 i5__i8__i10__net25 vss 47.8576e-18
c30 i5__i8__i9__net22 vss 46.2729e-18
c31 i5__i8__i9__net23 vss 114.453e-21
c32 i5__i8__i9__net24 vss 50.2132e-18
c33 i5__i8__i9__net21 vss 114.718e-21
c34 i5__i8__i9__net25 vss 49.2786e-18
c35 i5__i8__i8__net2 vss 97.9536e-18
c36 i5__i8__i8__net1 vss 29.6683e-18
c37 i5__i7__y1out vss 112.449e-18
c38 i5__i7__x1out vss 110.574e-18
c39 i5__i7__xor1 vss 36.6535e-18
c40 i5__i7__y0out vss 109.724e-18
c41 i5__i7__x0out vss 110.227e-18
c42 i5__i7__xor0 vss 32.0032e-18
c43 i5__i7__y2out vss 31.4762e-18
c44 i5__i7__x2out vss 35.4091e-18
c45 i5__i7__xor2 vss 38.7719e-18
c46 i5__i7__y3out vss 31.3786e-18
c47 i5__i7__x3out vss 35.2645e-18
c48 i5__i7__xor3 vss 31.0412e-18
c49 i5__i7__net44 vss 35.739e-18
c50 i5__i7__net47 vss 31.6164e-18
c51 i5__i7__net46 vss 35.3892e-18
c52 i5__i7__net50 vss 32.117e-18
c53 i5__i7__net51 vss 37.9289e-18
c54 i5__i7__i1__net1 vss 20.743e-18
c55 i5__i7__i1__i2__net25 vss 52.4503e-18
c56 i5__i7__i1__i2__net24 vss 68.8373e-18
c57 i5__i7__i1__i2__net22 vss 26.0494e-18
c58 i5__i7__i1__i2__net23 vss 52.4491e-18
c59 i5__i7__i1__i2__net21 vss 66.8397e-18
c60 i5__i7__i1__i1__net25 vss 53.039e-18
c61 i5__i7__i1__i1__net24 vss 69.4201e-18
c62 i5__i7__i1__i1__net22 vss 25.3565e-18
c63 i5__i7__i1__i1__net23 vss 52.829e-18
c64 i5__i7__i1__i1__net21 vss 67.0466e-18
c65 i5__i7__i1__i0__net25 vss 52.9076e-18
c66 i5__i7__i1__i0__net24 vss 69.3193e-18
c67 i5__i7__i1__i0__net22 vss 25.4692e-18
c68 i5__i7__i1__i0__net23 vss 52.8369e-18
c69 i5__i7__i1__i0__net21 vss 68.5264e-18
c70 i5__i7__i1__i3__net25 vss 52.9843e-18
c71 i5__i7__i1__i3__net24 vss 69.7241e-18
c72 i5__i7__i1__i3__net22 vss 24.8145e-18
c73 i5__i7__i1__i3__net23 vss 54.7415e-18
c74 i5__i7__i1__i3__net21 vss 69.4219e-18
c75 i5__i7__i0__net1 vss 20.3333e-18
c76 i5__i7__i0__i2__net25 vss 52.6152e-18
c77 i5__i7__i0__i2__net24 vss 67.6491e-18
c78 i5__i7__i0__i2__net22 vss 23.755e-18
c79 i5__i7__i0__i2__net23 vss 52.8103e-18
c80 i5__i7__i0__i2__net21 vss 65.7612e-18
c81 i5__i7__i0__i1__net25 vss 53.1755e-18
c82 i5__i7__i0__i1__net24 vss 69.6505e-18
c83 i5__i7__i0__i1__net22 vss 24.6127e-18
c84 i5__i7__i0__i1__net23 vss 52.8247e-18
c85 i5__i7__i0__i1__net21 vss 64.8674e-18
c86 i5__i7__i0__i0__net25 vss 53.0821e-18
c87 i5__i7__i0__i0__net24 vss 69.6832e-18
c88 i5__i7__i0__i0__net22 vss 25.1108e-18
c89 i5__i7__i0__i0__net23 vss 52.921e-18
c90 i5__i7__i0__i0__net21 vss 66.3571e-18
c91 i5__i7__i0__i3__net25 vss 52.7892e-18
c92 i5__i7__i0__i3__net24 vss 72.3861e-18
c93 i5__i7__i0__i3__net22 vss 23.7893e-18
c94 i5__i7__i0__i3__net23 vss 55.9801e-18
c95 i5__i7__i0__i3__net21 vss 69.8133e-18
c96 i5__i7__i5__net1 vss 38.1505e-18
c97 i5__i7__i6__net1 vss 38.3922e-18
c98 i5__i7__i4__net1 vss 36.6927e-18
c99 i5__i7__i7__net3 vss 33.6965e-18
c100 i5__i7__i7__net1 vss 30.2065e-18
c101 i5__i7__i7__net2 vss 37.1e-18
c102 i5__i7__i7__i1__net1 vss 25.6721e-18
c103 i5__i7__i7__i0__net1 vss 26.2625e-18
c104 i5__i7__i7__i4__net2 vss 92.9707e-18
c105 i5__i7__i7__i4__net3 vss 84.9499e-18
c106 i5__i7__i7__i4__net4 vss 64.3116e-18
c107 i5__i7__i7__i4__net1 vss 69.4946e-18
c108 i5__i7__i9__net1 vss 25.6935e-18
c109 i5__i7__i8__net1 vss 26.5267e-18
c110 i5__i7__i2__net1 vss 25.796e-18
c111 i5__i7__i3__net1 vss 26.6186e-18
c112 i5__i9__net21 vss 55.5512e-18
c113 i5__i6__net30 vss 45.0878e-18
c114 i5__i6__net32 vss 74.2349e-18
c115 i5__i6__net33 vss 45.8516e-18
c116 i5__i6__net34 vss 73.8641e-18
c117 i5__i6__net35 vss 43.8576e-18
c118 i5__i6__net31 vss 32.9406e-18
c119 i5__i6__i5__net22 vss 43.872e-18
c120 i5__i6__i5__net23 vss 12.2584e-21
c121 i5__i6__i5__net24 vss 50.8661e-18
c122 i5__i6__i5__net21 vss 545.681e-21
c123 i5__i6__i5__net25 vss 56.6281e-18
c124 i5__i6__i4__net22 vss 45.2369e-18
c125 i5__i6__i4__net24 vss 50.094e-18
c126 i5__i6__i4__net21 vss 151.115e-21
c127 i5__i6__i4__net25 vss 55.6154e-18
c128 i5__i6__i2__net22 vss 44.6603e-18
c129 i5__i6__i2__net23 vss 409.378e-21
c130 i5__i6__i2__net24 vss 51.3243e-18
c131 i5__i6__i2__net21 vss 517.697e-21
c132 i5__i6__i2__net25 vss 56.4789e-18
c133 i5__i6__i8__net4 vss 20.5012e-18
c134 i5__i6__i7__net4 vss 20.3745e-18
c135 i5__i6__i6__net4 vss 20.2934e-18
c136 i4__net1 vss 48.7633e-18
c137 i1__net4 vss 44.724e-18
c138 i1__net3 vss 328.221e-18
c139 i1__net2 vss 21.3653e-18
c140 i1__i14__net1 vss 253.247e-18
c141 i1__i11__outinv vss 30.7981e-18
c142 i1__i13__net1 vss 143.998e-18
c143 i1__i12__net1 vss 37.9621e-18
c144 n52__i1__net3 vss 158.139e-18
c145 n48__i1__net3 vss 150.164e-18
c146 n44__i1__net3 vss 153.783e-18
c147 n40__i1__net3 vss 152.587e-18
c148 n36__i1__net3 vss 155.347e-18
c149 n32__i1__net3 vss 159.676e-18
c150 n121__i1__i13__net1 vss 170.228e-18
c151 n4__i1__i11__outinv vss 28.6401e-18
c152 n97__i1__i13__net1 vss 155.056e-18
c153 n2__i1__i11__outinv vss 33.8022e-18
c154 n89__i1__i13__net1 vss 155.219e-18
c155 n81__i1__i13__net1 vss 155.16e-18
c156 n77__i1__i13__net1 vss 160.392e-18
c157 n65__i1__i13__net1 vss 161.912e-18
c158 n12__i1__net4 vss 35.5475e-18
c159 n57__i1__i13__net1 vss 162.881e-18
c160 n10__i1__net4 vss 41.4706e-18
c161 n53__i1__i13__net1 vss 160.509e-18
c162 n49__i1__i13__net1 vss 159.569e-18
c163 n45__i1__i13__net1 vss 157.759e-18
c164 n7__i1__net4 vss 72.1778e-18
c165 n41__i1__i13__net1 vss 158.016e-18
c166 n3__i1__net4 vss 63.6028e-18
c167 n37__i1__i13__net1 vss 159.314e-18
c168 n33__i1__i13__net1 vss 162.074e-18
c169 n29__i1__i13__net1 vss 158.213e-18
c170 n27__i1__i12__net1 vss 70.5406e-18
c171 n25__i1__i13__net1 vss 156.423e-18
c172 n23__i1__i12__net1 vss 54.7278e-18
c173 n21__i1__i13__net1 vss 154.49e-18
c174 n19__i1__i12__net1 vss 51.553e-18
c175 n17__i1__i13__net1 vss 155.168e-18
c176 n15__i1__i12__net1 vss 56.5805e-18
c177 n13__i1__i13__net1 vss 158.131e-18
c178 n11__i1__i12__net1 vss 57.8831e-18
c179 n9__i1__i13__net1 vss 161.712e-18
c180 n7__i1__i12__net1 vss 59.1366e-18
c181 n5__i1__i13__net1 vss 157.504e-18
c182 n3__i1__i12__net1 vss 48.0764e-18
c183 n183__i1__net2 vss 352.895e-18
c184 n155__i1__net2 vss 323.853e-18
c185 n147__i1__net2 vss 381.92e-18
c186 n139__i1__net2 vss 331.981e-18
c187 n135__i1__net2 vss 381.087e-18
c188 n123__i1__net2 vss 329.729e-18
c189 n115__i1__net2 vss 381.892e-18
c190 n107__i1__net2 vss 317.398e-18
c191 n103__i1__net2 vss 381.629e-18
c192 n95__i1__net2 vss 321.107e-18
c193 n87__i1__net2 vss 380.448e-18
c194 n75__i1__net2 vss 330.592e-18
c195 n67__i1__net2 vss 382.398e-18
c196 n59__i1__net2 vss 327.498e-18
c197 n55__i1__net2 vss 381.914e-18
c198 n51__i1__net2 vss 333.599e-18
c199 n47__i1__net2 vss 341.747e-18
c200 n43__i1__net2 vss 377.406e-18
c201 n39__i1__net2 vss 331.419e-18
c202 n35__i1__net2 vss 375.267e-18
c203 n31__i1__net2 vss 324.663e-18
c204 n27__i1__net2 vss 388.729e-18
c205 n23__i1__net2 vss 335.001e-18
c206 n19__i1__net2 vss 390.583e-18
c207 n15__i1__net2 vss 339.968e-18
c208 n12__i1__net2 vss 377.466e-18
c209 n7__i1__net2 vss 332.545e-18
c210 n4__i1__net2 vss 313.802e-18
c211 n715__i1__i14__net1 vss 408.465e-18
c212 n707__i1__i14__net1 vss 327.842e-18
c213 n703__i1__i14__net1 vss 385.159e-18
c214 n691__i1__i14__net1 vss 374.609e-18
c215 n687__i1__i14__net1 vss 364.879e-18
c216 n675__i1__i14__net1 vss 369.855e-18
c217 n671__i1__i14__net1 vss 366.614e-18
c218 n659__i1__i14__net1 vss 325.956e-18
c219 n651__i1__i14__net1 vss 380.004e-18
c220 n647__i1__i14__net1 vss 326.046e-18
c221 n639__i1__i14__net1 vss 381.287e-18
c222 n631__i1__i14__net1 vss 370.437e-18
c223 n619__i1__i14__net1 vss 365.119e-18
c224 n611__i1__i14__net1 vss 374.617e-18
c225 n607__i1__i14__net1 vss 365.9e-18
c226 n595__i1__i14__net1 vss 363.932e-18
c227 n591__i1__i14__net1 vss 364.177e-18
c228 n579__i1__i14__net1 vss 348.396e-18
c229 n571__i1__i14__net1 vss 366.137e-18
c230 n563__i1__i14__net1 vss 346.939e-18
c231 n555__i1__i14__net1 vss 325.803e-18
c232 n547__i1__i14__net1 vss 367.345e-18
c233 n543__i1__i14__net1 vss 326.122e-18
c234 n531__i1__i14__net1 vss 360.958e-18
c235 n527__i1__i14__net1 vss 357.456e-18
c236 n515__i1__i14__net1 vss 348.16e-18
c237 n507__i1__i14__net1 vss 367.523e-18
c238 n499__i1__i14__net1 vss 352.754e-18
c239 n495__i1__i14__net1 vss 325.711e-18
c240 n483__i1__i14__net1 vss 368.3e-18
c241 n479__i1__i14__net1 vss 366.838e-18
c242 n467__i1__i14__net1 vss 355.115e-18
c243 n459__i1__i14__net1 vss 374.814e-18
c244 n451__i1__i14__net1 vss 381.464e-18
c245 n443__i1__i14__net1 vss 335.257e-18
c246 n435__i1__i14__net1 vss 390.459e-18
c247 n427__i1__i14__net1 vss 340.02e-18
c248 n424__i1__i14__net1 vss 376.955e-18
c249 n415__i1__i14__net1 vss 380.042e-18
c250 n408__i1__i14__net1 vss 362.048e-18
c251 n395__i1__i14__net1 vss 373.404e-18
c252 n392__i1__i14__net1 vss 379.802e-18
c253 n381__i1__i14__net1 vss 333.997e-18
c254 n376__i1__i14__net1 vss 389.911e-18
c255 n363__i1__i14__net1 vss 335.257e-18
c256 n360__i1__i14__net1 vss 378.059e-18
c257 n347__i1__i14__net1 vss 381.223e-18
c258 n344__i1__i14__net1 vss 328.139e-18
c259 n335__i1__i14__net1 vss 381.913e-18
c260 n328__i1__i14__net1 vss 326.218e-18
c261 n315__i1__i14__net1 vss 366.082e-18
c262 n308__i1__i14__net1 vss 366.72e-18
c263 n303__i1__i14__net1 vss 364.58e-18
c264 n295__i1__i14__net1 vss 372.529e-18
c265 n287__i1__i14__net1 vss 381.359e-18
c266 n275__i1__i14__net1 vss 324.756e-18
c267 n271__i1__i14__net1 vss 382.397e-18
c268 n259__i1__i14__net1 vss 325.902e-18
c269 n255__i1__i14__net1 vss 381.93e-18
c270 n243__i1__i14__net1 vss 320.624e-18
c271 n239__i1__i14__net1 vss 379.855e-18
c272 n227__i1__i14__net1 vss 335.271e-18
c273 n219__i1__i14__net1 vss 380.771e-18
c274 n211__i1__i14__net1 vss 326.038e-18
c275 n203__i1__i14__net1 vss 380.601e-18
c276 n199__i1__i14__net1 vss 317.182e-18
c277 n187__i1__i14__net1 vss 381.593e-18
c278 n179__i1__i14__net1 vss 323.008e-18
c279 n175__i1__i14__net1 vss 381.744e-18
c280 n163__i1__i14__net1 vss 332.037e-18
c281 n159__i1__i14__net1 vss 382.355e-18
c282 n147__i1__i14__net1 vss 326.973e-18
c283 n143__i1__i14__net1 vss 378.956e-18
c284 n133__i1__i14__net1 vss 328.604e-18
c285 n127__i1__i14__net1 vss 338.283e-18
c286 n115__i1__i14__net1 vss 381.767e-18
c287 n107__i1__i14__net1 vss 331.246e-18
c288 n99__i1__i14__net1 vss 373.449e-18
c289 n91__i1__i14__net1 vss 322.961e-18
c290 n83__i1__i14__net1 vss 378.33e-18
c291 n79__i1__i14__net1 vss 332.063e-18
c292 n68__i1__i14__net1 vss 373.509e-18
c293 n59__i1__i14__net1 vss 337.286e-18
c294 n56__i1__i14__net1 vss 368.802e-18
c295 n51__i1__i14__net1 vss 328.118e-18
c296 n48__i1__i14__net1 vss 369.085e-18
c297 n43__i1__i14__net1 vss 319.138e-18
c298 n40__i1__i14__net1 vss 375.621e-18
c299 n35__i1__i14__net1 vss 358.024e-18
c300 n32__i1__i14__net1 vss 370.035e-18
c301 n27__i1__i14__net1 vss 376.847e-18
c302 n24__i1__i14__net1 vss 323.047e-18
c303 n19__i1__i14__net1 vss 377.288e-18
c304 n15__i1__i14__net1 vss 322.783e-18
c305 n11__i1__i14__net1 vss 376.905e-18
c306 n7__i1__i14__net1 vss 322.257e-18
c307 n3__i1__i14__net1 vss 389.988e-18
c308 n1__piso_out vss 26.7227e-18
c309 n9__piso_out vss 18.2667e-18
c310 n11__piso_out vss 16.8818e-18
c311 n30__i5__i8__net2 vss 59.4721e-18
c312 n13__piso_out vss 19.9658e-18
c313 n85__i5__clk4 vss 44.1063e-18
c314 n5__i4__net1 vss 28.8369e-18
c315 n76__i5__clk4 vss 21.1415e-18
c316 n80__i5__clk4 vss 13.8292e-18
c317 n78__i5__clk4 vss 22.4931e-18
c318 n15__i5__i8__net1 vss 42.941e-18
c319 n38__i5__i6__net31 vss 37.7617e-18
c320 n16__i5__i8__net1 vss 39.2935e-18
c321 n39__i5__i6__net31 vss 39.3666e-18
c322 n6__i5__i8__i10__net22 vss 21.4505e-18
c323 n6__i5__i6__i5__net22 vss 21.4617e-18
c324 n10__i5__i8__net2 vss 34.7224e-18
c325 n53__i5__clk_buf vss 33.0912e-18
c326 n11__i5__i8__net2 vss 47.9708e-18
c327 n54__i5__clk_buf vss 46.398e-18
c328 n6__i5__i8__net5 vss 26.5875e-18
c329 n6__i5__i6__net35 vss 26.0227e-18
c330 n32__shift vss 20.9533e-18
c331 n5__i5__i8__net2 vss 13.6331e-18
c332 n3__i5__i8__net2 vss 23.0381e-18
c333 n23__shift vss 24.8172e-18
c334 n5__i5__i8__net4 vss 38.2698e-18
c335 n6__i5__i8__net4 vss 39.3212e-18
c336 n6__i5__i8__i9__net22 vss 26.3939e-18
c337 n26__i5__i6__net31 vss 42.7307e-18
c338 n27__i5__i6__net31 vss 39.3948e-18
c339 n32__i5__clk_buf vss 34.9387e-18
c340 n6__i5__i6__i4__net22 vss 21.3975e-18
c341 n33__i5__clk_buf vss 45.8903e-18
c342 n6__i5__i8__net1 vss 25.1451e-18
c343 n29__i5__clk_buf vss 33.4213e-18
c344 n30__i5__clk_buf vss 46.2561e-18
c345 n18__i5__clk_buf vss 22.3429e-18
c346 n6__i5__i6__net33 vss 26.7171e-18
c347 n22__i5__clk_buf vss 12.3438e-18
c348 n20__i5__clk_buf vss 23.9245e-18
c349 n19__shift vss 20.6997e-18
c350 n15__i5__i9__net21 vss 25.0787e-18
c351 n11__i5__i9__net21 vss 15.8183e-18
c352 n7__i5__i9__net21 vss 17.3987e-18
c353 n2__i5__i9__net21 vss 16.3605e-18
c354 n10__shift vss 25.1097e-18
c355 n1__clk_out vss 42.4576e-18
c356 n5__clk_out vss 30.5068e-18
c357 n5__i5__i6__net31 vss 42.025e-18
c358 n6__i5__i6__net31 vss 39.262e-18
c359 n6__i5__i6__i2__net22 vss 21.0404e-18
c360 n20__i5__i7__net44 vss 37.4711e-18
c361 n10__i5__clk_buf vss 32.3112e-18
c362 n11__i5__clk_buf vss 45.6782e-18
c363 n15__i5__i7__i7__net1 vss 33.058e-18
c364 n8__i5__i7__net46 vss 33.8747e-18
c365 n6__i5__i6__net30 vss 26.0789e-18
c366 n6__shift vss 21.6073e-18
c367 n6__i5__i7__i7__net1 vss 30.8571e-18
c368 n1__shift vss 21.831e-18
c369 n4__i5__i7__i7__net1 vss 25.119e-18
c370 n5__i5__clk_buf vss 12.2719e-18
c371 n3__i5__clk_buf vss 22.9747e-18
c372 n6__i5__i7__net51 vss 22.7533e-18
c373 n4__i5__i7__net47 vss 24.5417e-18
c374 n13__i5__i7__xor2 vss 24.0287e-18
c375 n13__i5__i7__xor1 vss 23.5132e-18
c376 n4__i5__i7__y3out vss 25.1958e-18
c377 n11__i5__i7__y0out vss 25.1241e-18
c378 n8__i5__i7__x0out vss 36.3348e-18
c379 n8__i5__i7__y0out vss 29.7652e-18
c380 n11__i5__i7__y2out vss 25.1463e-18
c381 n11__i5__i7__y1out vss 24.9747e-18
c382 n8__i5__i7__x1out vss 36.3497e-18
c383 n8__i5__i7__y1out vss 29.8286e-18
c384 n25__i5__i7__i1__net1 vss 24.5033e-18
c385 n25__i5__i7__i0__net1 vss 24.4399e-18
c386 n48__i5__clk4 vss 23.2629e-18
c387 n46__i5__clk4 vss 23.1862e-18
c388 n1__y3 vss 25.1181e-18
c389 n1__x3 vss 24.8813e-18
c390 n18__i5__i7__i1__net1 vss 24.1794e-18
c391 n18__i5__i7__i0__net1 vss 24.2565e-18
c392 n38__i5__clk4 vss 23.1562e-18
c393 n36__i5__clk4 vss 23.1472e-18
c394 n1__y2 vss 25.6599e-18
c395 n1__x2 vss 26.1018e-18
c396 n11__i5__i7__i1__net1 vss 24.338e-18
c397 n11__i5__i7__i0__net1 vss 24.8435e-18
c398 n17__i5__clk4 vss 23.1948e-18
c399 n15__i5__clk4 vss 23.195e-18
c400 n1__y1 vss 25.4452e-18
c401 n1__x1 vss 25.4651e-18
c402 n3__i5__i7__i1__net1 vss 24.3579e-18
c403 n3__i5__i7__i0__net1 vss 23.9537e-18
c404 n9__i5__clk4 vss 23.3868e-18
c405 n7__i5__clk4 vss 23.3756e-18
c406 n1__y0 vss 23.16e-18
c407 n1__x0 vss 22.3701e-18
c408 n4__i5__clk4 vss 38.9389e-18
c409 n50__i1__net3 vss 115.222e-18
c410 n46__i1__net3 vss 111.975e-18
c411 n42__i1__net3 vss 115.631e-18
c412 n38__i1__net3 vss 115.868e-18
c413 n34__i1__net3 vss 116.374e-18
c414 n30__i1__net3 vss 120.602e-18
c415 n124__i1__i13__net1 vss 115.399e-18
c416 n14__piso_outinv vss 54.8224e-18
c417 n99__i1__i13__net1 vss 109.821e-18
c418 n12__piso_outinv vss 43.5465e-18
c419 n92__i1__i13__net1 vss 109.901e-18
c420 n10__piso_outinv vss 49.0018e-18
c421 n83__i1__i13__net1 vss 111.357e-18
c422 n80__i1__i13__net1 vss 109.425e-18
c423 n27__piso_out vss 51.5202e-18
c424 n67__i1__i13__net1 vss 108.608e-18
c425 n25__piso_out vss 41.7526e-18
c426 n60__i1__i13__net1 vss 118.298e-18
c427 n22__piso_out vss 47.3372e-18
c428 n55__i1__i13__net1 vss 117.176e-18
c429 n52__i1__i13__net1 vss 115.472e-18
c430 n47__i1__i13__net1 vss 116.774e-18
c431 n5__i1__net4 vss 51.3636e-18
c432 n44__i1__i13__net1 vss 117.029e-18
c433 n39__i1__i13__net1 vss 119.338e-18
c434 n36__i1__i13__net1 vss 117.591e-18
c435 n31__i1__i13__net1 vss 112.996e-18
c436 n25__i1__i12__net1 vss 48.9593e-18
c437 n28__i1__i13__net1 vss 110.908e-18
c438 n21__i1__i12__net1 vss 39.9993e-18
c439 n23__i1__i13__net1 vss 113.49e-18
c440 n17__i1__i12__net1 vss 37.904e-18
c441 n19__i1__i13__net1 vss 111.412e-18
c442 n13__i1__i12__net1 vss 41.428e-18
c443 n15__i1__i13__net1 vss 110.39e-18
c444 n9__i1__i12__net1 vss 41.4539e-18
c445 n11__i1__i13__net1 vss 114.351e-18
c446 n5__i1__i12__net1 vss 39.2286e-18
c447 n7__i1__i13__net1 vss 116.705e-18
c448 n3__i1__i13__net1 vss 108.63e-18
c449 n181__i1__net2 vss 246.542e-18
c450 n153__i1__net2 vss 214.852e-18
c451 n145__i1__net2 vss 253.46e-18
c452 n137__i1__net2 vss 213.635e-18
c453 n133__i1__net2 vss 251.669e-18
c454 n121__i1__net2 vss 213.527e-18
c455 n113__i1__net2 vss 254.42e-18
c456 n105__i1__net2 vss 214.979e-18
c457 n101__i1__net2 vss 254.635e-18
c458 n93__i1__net2 vss 214.589e-18
c459 n85__i1__net2 vss 254.597e-18
c460 n73__i1__net2 vss 214.5e-18
c461 n65__i1__net2 vss 254.152e-18
c462 n57__i1__net2 vss 215.176e-18
c463 n53__i1__net2 vss 252.879e-18
c464 n49__i1__net2 vss 225.839e-18
c465 n45__i1__net2 vss 255.118e-18
c466 n41__i1__net2 vss 215.943e-18
c467 n37__i1__net2 vss 256.935e-18
c468 n33__i1__net2 vss 216.028e-18
c469 n29__i1__net2 vss 256.69e-18
c470 n25__i1__net2 vss 216.139e-18
c471 n21__i1__net2 vss 256.979e-18
c472 n17__i1__net2 vss 215.55e-18
c473 n13__i1__net2 vss 255.009e-18
c474 n10__i1__net2 vss 213.983e-18
c475 n5__i1__net2 vss 254.563e-18
c476 n2__i1__net2 vss 234.643e-18
c477 n713__i1__i14__net1 vss 235.719e-18
c478 n705__i1__i14__net1 vss 212.4e-18
c479 n701__i1__i14__net1 vss 250.614e-18
c480 n689__i1__i14__net1 vss 217.52e-18
c481 n685__i1__i14__net1 vss 252.011e-18
c482 n673__i1__i14__net1 vss 215.21e-18
c483 n669__i1__i14__net1 vss 255.047e-18
c484 n657__i1__i14__net1 vss 210.768e-18
c485 n649__i1__i14__net1 vss 252.637e-18
c486 n645__i1__i14__net1 vss 212.879e-18
c487 n637__i1__i14__net1 vss 252.639e-18
c488 n629__i1__i14__net1 vss 215.968e-18
c489 n617__i1__i14__net1 vss 252.204e-18
c490 n609__i1__i14__net1 vss 211.814e-18
c491 n605__i1__i14__net1 vss 253.201e-18
c492 n593__i1__i14__net1 vss 220.593e-18
c493 n589__i1__i14__net1 vss 255.27e-18
c494 n577__i1__i14__net1 vss 214.992e-18
c495 n569__i1__i14__net1 vss 254.332e-18
c496 n561__i1__i14__net1 vss 216.707e-18
c497 n553__i1__i14__net1 vss 254.675e-18
c498 n545__i1__i14__net1 vss 214.692e-18
c499 n541__i1__i14__net1 vss 254.061e-18
c500 n529__i1__i14__net1 vss 210.034e-18
c501 n525__i1__i14__net1 vss 247.797e-18
c502 n513__i1__i14__net1 vss 212.952e-18
c503 n505__i1__i14__net1 vss 255.067e-18
c504 n497__i1__i14__net1 vss 215.112e-18
c505 n493__i1__i14__net1 vss 227.663e-18
c506 n481__i1__i14__net1 vss 247.767e-18
c507 n477__i1__i14__net1 vss 218.632e-18
c508 n465__i1__i14__net1 vss 252.647e-18
c509 n457__i1__i14__net1 vss 219.601e-18
c510 n449__i1__i14__net1 vss 248.727e-18
c511 n441__i1__i14__net1 vss 217.718e-18
c512 n433__i1__i14__net1 vss 245.526e-18
c513 n425__i1__i14__net1 vss 217.96e-18
c514 n422__i1__i14__net1 vss 247.812e-18
c515 n413__i1__i14__net1 vss 218.259e-18
c516 n406__i1__i14__net1 vss 252.338e-18
c517 n393__i1__i14__net1 vss 217.566e-18
c518 n390__i1__i14__net1 vss 253.491e-18
c519 n379__i1__i14__net1 vss 219.359e-18
c520 n374__i1__i14__net1 vss 247.868e-18
c521 n361__i1__i14__net1 vss 248.521e-18
c522 n358__i1__i14__net1 vss 241.784e-18
c523 n345__i1__i14__net1 vss 243.174e-18
c524 n342__i1__i14__net1 vss 242.496e-18
c525 n333__i1__i14__net1 vss 243.982e-18
c526 n326__i1__i14__net1 vss 246.723e-18
c527 n313__i1__i14__net1 vss 246.5e-18
c528 n306__i1__i14__net1 vss 247.806e-18
c529 n301__i1__i14__net1 vss 244.966e-18
c530 n293__i1__i14__net1 vss 243.461e-18
c531 n285__i1__i14__net1 vss 247.292e-18
c532 n273__i1__i14__net1 vss 240.457e-18
c533 n269__i1__i14__net1 vss 244.018e-18
c534 n257__i1__i14__net1 vss 212.871e-18
c535 n253__i1__i14__net1 vss 216.758e-18
c536 n241__i1__i14__net1 vss 244.285e-18
c537 n237__i1__i14__net1 vss 241.955e-18
c538 n225__i1__i14__net1 vss 244.694e-18
c539 n217__i1__i14__net1 vss 254.133e-18
c540 n209__i1__i14__net1 vss 216.169e-18
c541 n201__i1__i14__net1 vss 245.793e-18
c542 n197__i1__i14__net1 vss 245.137e-18
c543 n185__i1__i14__net1 vss 242.463e-18
c544 n177__i1__i14__net1 vss 242.012e-18
c545 n173__i1__i14__net1 vss 242.07e-18
c546 n161__i1__i14__net1 vss 245.279e-18
c547 n157__i1__i14__net1 vss 245.581e-18
c548 n145__i1__i14__net1 vss 245.25e-18
c549 n141__i1__i14__net1 vss 244.145e-18
c550 n131__i1__i14__net1 vss 238.062e-18
c551 n125__i1__i14__net1 vss 250.704e-18
c552 n113__i1__i14__net1 vss 219.351e-18
c553 n105__i1__i14__net1 vss 253.797e-18
c554 n97__i1__i14__net1 vss 212.45e-18
c555 n89__i1__i14__net1 vss 251.703e-18
c556 n81__i1__i14__net1 vss 211.647e-18
c557 n77__i1__i14__net1 vss 251.771e-18
c558 n66__i1__i14__net1 vss 213.686e-18
c559 n57__i1__i14__net1 vss 251.061e-18
c560 n54__i1__i14__net1 vss 212.668e-18
c561 n49__i1__i14__net1 vss 251.075e-18
c562 n46__i1__i14__net1 vss 212.93e-18
c563 n41__i1__i14__net1 vss 245.828e-18
c564 n38__i1__i14__net1 vss 245.841e-18
c565 n33__i1__i14__net1 vss 213.32e-18
c566 n30__i1__i14__net1 vss 250.736e-18
c567 n25__i1__i14__net1 vss 220.506e-18
c568 n22__i1__i14__net1 vss 246.877e-18
c569 n17__i1__i14__net1 vss 219.81e-18
c570 n13__i1__i14__net1 vss 246.494e-18
c571 n9__i1__i14__net1 vss 219.607e-18
c572 n5__i1__i14__net1 vss 250.341e-18
c573 n3__i5__i8__i8__net1 vss 21.163e-18
c574 n7__piso_out vss 25.7115e-18
c575 n8__piso_out vss 15.4354e-18
c576 n10__piso_out vss 14.4048e-18
c577 n31__i5__i8__net2 vss 32.0303e-18
c578 n12__piso_out vss 18.0786e-18
c579 n88__i5__clk4 vss 31.0643e-18
c580 n2__i4__net1 vss 36.7807e-18
c581 n3__i4__net1 vss 24.2782e-18
c582 n84__i5__clk4 vss 20.3975e-18
c583 n83__i5__clk4 vss 10.7425e-18
c584 n81__i5__clk4 vss 18.5162e-18
c585 n3__bufin vss 27.8625e-18
c586 n60__reset vss 35.8555e-18
c587 n56__reset vss 40.6752e-18
c588 n63__reset vss 24.6886e-18
c589 n59__reset vss 24.9032e-18
c590 n13__i5__i8__net2 vss 28.7762e-18
c591 n60__i5__clk_buf vss 31.516e-18
c592 n14__i5__i8__net2 vss 30.0238e-18
c593 n61__i5__clk_buf vss 29.9527e-18
c594 n7__i5__i8__i10__net22 vss 34.7342e-18
c595 n7__i5__i6__i5__net22 vss 37.9935e-18
c596 n5__i5__i8__i10__net22 vss 17.0714e-18
c597 n5__i5__i6__i5__net22 vss 20.3195e-18
c598 n11__i5__i8__net1 vss 29.3311e-18
c599 n32__i5__i6__net31 vss 32.0883e-18
c600 n14__i5__i8__net1 vss 21.6391e-18
c601 n35__i5__i6__net31 vss 25.0504e-18
c602 n7__i5__i8__net5 vss 30.9425e-18
c603 n7__i5__i6__net35 vss 34.508e-18
c604 n5__i5__i8__net5 vss 18.7965e-18
c605 n5__i5__i6__net35 vss 20.7705e-18
c606 n3__i5__i6__i8__net4 vss 18.2633e-18
c607 n9__i5__i8__net2 vss 20.4417e-18
c608 n8__i5__i8__net2 vss 11.5006e-18
c609 n6__i5__i8__net2 vss 19.1201e-18
c610 n30__shift vss 17.0768e-18
c611 n47__reset vss 37.0404e-18
c612 n25__shift vss 19.3425e-18
c613 n50__reset vss 25.3454e-18
c614 n43__reset vss 38.9395e-18
c615 n40__i5__clk_buf vss 28.1267e-18
c616 n46__reset vss 26.3176e-18
c617 n41__i5__clk_buf vss 29.761e-18
c618 n7__i5__i8__i9__net22 vss 35.0654e-18
c619 n5__i5__i8__i9__net22 vss 17.3378e-18
c620 n37__i5__clk_buf vss 32.13e-18
c621 n38__i5__clk_buf vss 30.6005e-18
c622 n7__i5__i6__i4__net22 vss 38.6748e-18
c623 n5__i5__i6__i4__net22 vss 19.2078e-18
c624 n4__i5__i8__net4 vss 22.1942e-18
c625 n7__i5__i8__net1 vss 32.2593e-18
c626 n5__i5__i8__net1 vss 19.6352e-18
c627 n18__i5__i6__net31 vss 32.2446e-18
c628 n21__i5__i6__net31 vss 25.1962e-18
c629 n7__i5__i6__net33 vss 34.898e-18
c630 n26__i5__clk_buf vss 23.2231e-18
c631 n5__i5__i6__net33 vss 20.7062e-18
c632 n25__i5__clk_buf vss 11.9189e-18
c633 n23__i5__clk_buf vss 21.3603e-18
c634 n3__i5__i6__i7__net4 vss 18.259e-18
c635 n17__i5__i9__net21 vss 18.6918e-18
c636 n17__shift vss 16.7727e-18
c637 n13__i5__i9__net21 vss 11.8158e-18
c638 n9__i5__i9__net21 vss 11.5455e-18
c639 n4__i5__i9__net21 vss 11.2901e-18
c640 n12__shift vss 18.2764e-18
c641 n2__clk_out vss 33.9391e-18
c642 n36__reset vss 38.5699e-18
c643 n3__clk_out vss 27.1062e-18
c644 n39__reset vss 25.6825e-18
c645 n13__i5__clk_buf vss 32.8215e-18
c646 n3__i5__i7__i7__net3 vss 27.0652e-18
c647 n14__i5__clk_buf vss 30.8125e-18
c648 n7__i5__i6__i2__net22 vss 39.071e-18
c649 n5__i5__i6__i2__net22 vss 19.2323e-18
c650 n18__i5__i7__i7__net1 vss 34.2948e-18
c651 n4__i5__i6__net31 vss 26.0266e-18
c652 n11__i5__i7__net46 vss 31.1087e-18
c653 n7__i5__i6__net30 vss 35.6545e-18
c654 n3__i5__i7__i7__net2 vss 29.974e-18
c655 n5__i5__i6__net30 vss 22.9442e-18
c656 n10__i5__i7__net44 vss 33.2973e-18
c657 n3__i5__i6__i6__net4 vss 18.1908e-18
c658 n4__shift vss 16.7976e-18
c659 n8__i5__i7__i7__net1 vss 25.2953e-18
c660 n3__shift vss 21.7605e-18
c661 n9__i5__clk_buf vss 26.7412e-18
c662 n8__i5__clk_buf vss 11.9821e-18
c663 n6__i5__clk_buf vss 20.6542e-18
c664 n3__i5__i7__net46 vss 37.8029e-18
c665 n5__i5__i7__i6__net1 vss 22.4814e-18
c666 n3__i5__i7__i7__net1 vss 21.4782e-18
c667 n3__i5__i7__net50 vss 40.246e-18
c668 n5__i5__i7__net51 vss 44.1204e-18
c669 n4__i5__i7__i6__net1 vss 41.1803e-18
c670 n3__i5__i7__net44 vss 39.9371e-18
c671 n3__i5__i7__net47 vss 22.6606e-18
c672 n3__i5__i7__net51 vss 24.9199e-18
c673 n5__i5__i7__i5__net1 vss 26.6257e-18
c674 n5__i5__i7__i4__net1 vss 26.9883e-18
c675 n3__i5__i7__xor3 vss 40.7007e-18
c676 n3__i5__i7__xor0 vss 40.4519e-18
c677 n12__i5__i7__xor2 vss 44.0651e-18
c678 n12__i5__i7__xor1 vss 43.9981e-18
c679 n4__i5__i7__i5__net1 vss 40.3185e-18
c680 n4__i5__i7__i4__net1 vss 41.4641e-18
c681 n3__i5__i7__xor2 vss 24.5829e-18
c682 n3__i5__i7__xor1 vss 25.0611e-18
c683 n3__i5__i7__x3out vss 38.1161e-18
c684 n10__i5__i7__x0out vss 38.8061e-18
c685 n3__i5__i7__y3out vss 21.7735e-18
c686 n10__i5__i7__y0out vss 22.0844e-18
c687 n3__i5__i7__x2out vss 40.8198e-18
c688 n10__i5__i7__x1out vss 40.0662e-18
c689 n3__i5__i7__y2out vss 19.2462e-18
c690 n10__i5__i7__y1out vss 19.3684e-18
c691 n26__reset vss 44.092e-18
c692 n24__reset vss 38.6242e-18
c693 n56__i5__clk4 vss 19.6425e-18
c694 n54__i5__clk4 vss 19.625e-18
c695 n4__i5__i7__i1__i2__net22 vss 25.894e-18
c696 n4__i5__i7__i0__i2__net22 vss 25.3001e-18
c697 n21__i5__i7__i1__net1 vss 21.1737e-18
c698 n21__i5__i7__i0__net1 vss 20.2194e-18
c699 n4__y3 vss 21.3598e-18
c700 n4__x3 vss 20.8944e-18
c701 n18__reset vss 40.9131e-18
c702 n16__reset vss 39.6024e-18
c703 n42__i5__clk4 vss 19.6529e-18
c704 n40__i5__clk4 vss 19.625e-18
c705 n4__i5__i7__i1__i1__net22 vss 25.3231e-18
c706 n4__i5__i7__i0__i1__net22 vss 24.6199e-18
c707 n16__i5__i7__i1__net1 vss 20.7729e-18
c708 n16__i5__i7__i0__net1 vss 20.2016e-18
c709 n4__y2 vss 20.5686e-18
c710 n4__x2 vss 20.7647e-18
c711 n7__reset vss 40.5618e-18
c712 n5__reset vss 39.4079e-18
c713 n28__i5__clk4 vss 20.0093e-18
c714 n26__i5__clk4 vss 20.1075e-18
c715 n4__i5__i7__i1__i0__net22 vss 25.3243e-18
c716 n4__i5__i7__i0__i0__net22 vss 25.538e-18
c717 n5__i5__i7__i1__net1 vss 20.7671e-18
c718 n5__i5__i7__i0__net1 vss 20.3574e-18
c719 n4__y1 vss 21.0738e-18
c720 n4__x1 vss 20.7407e-18
c721 n3__reset vss 40.2492e-18
c722 n1__reset vss 39.7272e-18
c723 n13__i5__clk4 vss 19.9621e-18
c724 n11__i5__clk4 vss 20.196e-18
c725 n4__i5__i7__i1__i3__net22 vss 25.0841e-18
c726 n4__i5__i7__i0__i3__net22 vss 25.4662e-18
c727 n4__y0 vss 25.1646e-18
c728 n4__x0 vss 24.876e-18
c729 n6__i5__clk4 vss 23.3136e-18
c730 n3__i5__clk4 vss 21.9665e-18
c731 n51__i1__net3 vss 26.536e-18
c732 n53__i1__net3 vss 26.4559e-18
c733 n47__i1__net3 vss 15.7201e-18
c734 n49__i1__net3 vss 15.5385e-18
c735 n43__i1__net3 vss 15.3894e-18
c736 n45__i1__net3 vss 15.2623e-18
c737 n39__i1__net3 vss 15.5656e-18
c738 n41__i1__net3 vss 15.4611e-18
c739 n35__i1__net3 vss 15.6415e-18
c740 n37__i1__net3 vss 15.487e-18
c741 n31__i1__net3 vss 22.8853e-18
c742 n33__i1__net3 vss 23.4066e-18
c743 n123__i1__i13__net1 vss 23.3747e-18
c744 n122__i1__i13__net1 vss 22.6736e-18
c745 n13__piso_outinv vss 24.3135e-18
c746 n3__i1__i11__outinv vss 25.4005e-18
c747 n100__i1__i13__net1 vss 15.5433e-18
c748 n98__i1__i13__net1 vss 15.2136e-18
c749 n11__piso_outinv vss 15.4445e-18
c750 n91__i1__i13__net1 vss 15.1475e-18
c751 n90__i1__i13__net1 vss 15.0095e-18
c752 n9__piso_outinv vss 23.5308e-18
c753 n84__i1__i13__net1 vss 15.5433e-18
c754 n82__i1__i13__net1 vss 15.2136e-18
c755 n79__i1__i13__net1 vss 15.1475e-18
c756 n78__i1__i13__net1 vss 15.0008e-18
c757 n26__piso_out vss 118.678e-18
c758 n68__i1__i13__net1 vss 56.9807e-18
c759 n66__i1__i13__net1 vss 51.3221e-18
c760 n11__i1__net4 vss 29.2261e-18
c761 n24__piso_out vss 15.2651e-18
c762 n59__i1__i13__net1 vss 15.1475e-18
c763 n58__i1__i13__net1 vss 15.098e-18
c764 n9__i1__net4 vss 25.0313e-18
c765 n23__piso_out vss 18.988e-18
c766 n56__i1__i13__net1 vss 15.5433e-18
c767 n54__i1__i13__net1 vss 15.2882e-18
c768 n51__i1__i13__net1 vss 15.1475e-18
c769 n50__i1__i13__net1 vss 15.098e-18
c770 n48__i1__i13__net1 vss 15.5433e-18
c771 n46__i1__i13__net1 vss 15.2882e-18
c772 n6__i1__net4 vss 26.9849e-18
c773 n8__i1__net4 vss 23.7133e-18
c774 n43__i1__i13__net1 vss 15.1475e-18
c775 n42__i1__i13__net1 vss 15.098e-18
c776 n2__i1__net4 vss 27.2577e-18
c777 n4__i1__net4 vss 25.27e-18
c778 n40__i1__i13__net1 vss 15.5433e-18
c779 n38__i1__i13__net1 vss 15.2882e-18
c780 n35__i1__i13__net1 vss 15.1013e-18
c781 n34__i1__i13__net1 vss 15.0435e-18
c782 n32__i1__i13__net1 vss 79.2116e-18
c783 n30__i1__i13__net1 vss 51.1442e-18
c784 n26__i1__i12__net1 vss 78.9188e-18
c785 n28__i1__i12__net1 vss 64.0243e-18
c786 n27__i1__i13__net1 vss 79.5086e-18
c787 n26__i1__i13__net1 vss 49.9569e-18
c788 n22__i1__i12__net1 vss 16.2209e-18
c789 n24__i1__i12__net1 vss 16.0318e-18
c790 n24__i1__i13__net1 vss 15.7158e-18
c791 n22__i1__i13__net1 vss 15.4459e-18
c792 n18__i1__i12__net1 vss 16.2152e-18
c793 n20__i1__i12__net1 vss 16.0521e-18
c794 n20__i1__i13__net1 vss 80.2224e-18
c795 n18__i1__i13__net1 vss 50.3973e-18
c796 n14__i1__i12__net1 vss 16.2047e-18
c797 n16__i1__i12__net1 vss 16.0585e-18
c798 n16__i1__i13__net1 vss 15.3626e-18
c799 n14__i1__i13__net1 vss 15.4831e-18
c800 n10__i1__i12__net1 vss 16.1776e-18
c801 n12__i1__i12__net1 vss 16.0591e-18
c802 n12__i1__i13__net1 vss 15.201e-18
c803 n10__i1__i13__net1 vss 16.6193e-18
c804 n6__i1__i12__net1 vss 16.2953e-18
c805 n8__i1__i12__net1 vss 16.8155e-18
c806 n8__i1__i13__net1 vss 56.4077e-18
c807 n6__i1__i13__net1 vss 68.4581e-18
c808 n2__i1__i12__net1 vss 29.237e-18
c809 n4__i1__i12__net1 vss 28.5226e-18
c810 n4__i1__i13__net1 vss 15.5686e-18
c811 n2__i1__i13__net1 vss 23.5595e-18
c812 n182__i1__net2 vss 22.632e-18
c813 n184__i1__net2 vss 23.0008e-18
c814 n2__i5__i8__i8__net1 vss 82.8043e-18
c815 n154__i1__net2 vss 14.6021e-18
c816 n156__i1__net2 vss 14.6451e-18
c817 n146__i1__net2 vss 60.8182e-18
c818 n148__i1__net2 vss 54.4155e-18
c819 n32__i5__i8__net2 vss 29.685e-18
c820 n138__i1__net2 vss 14.5873e-18
c821 n140__i1__net2 vss 14.6155e-18
c822 n6__piso_out vss 147.34e-18
c823 n87__i5__clk4 vss 10.5356e-18
c824 n134__i1__net2 vss 14.5873e-18
c825 n136__i1__net2 vss 14.6155e-18
c826 n122__i1__net2 vss 14.5873e-18
c827 n124__i1__net2 vss 14.6155e-18
c828 n4__i4__net1 vss 71.9822e-18
c829 n114__i1__net2 vss 14.5873e-18
c830 n116__i1__net2 vss 14.6155e-18
c831 n79__i5__clk4 vss 80.94e-18
c832 n2__bufin vss 93.1178e-18
c833 n106__i1__net2 vss 14.4994e-18
c834 n108__i1__net2 vss 14.5279e-18
c835 n102__i1__net2 vss 14.3105e-18
c836 n104__i1__net2 vss 14.3389e-18
c837 n94__i1__net2 vss 37.9363e-18
c838 n96__i1__net2 vss 47.1499e-18
c839 n62__reset vss 31.7198e-18
c840 n58__reset vss 32.4296e-18
c841 n86__i1__net2 vss 14.3856e-18
c842 n88__i1__net2 vss 14.4137e-18
c843 n74__i1__net2 vss 14.1998e-18
c844 n76__i1__net2 vss 14.228e-18
c845 n17__i5__i8__net1 vss 22.7535e-18
c846 n15__i5__i8__net2 vss 26.5559e-18
c847 n40__i5__i6__net31 vss 23.9446e-18
c848 n62__i5__clk_buf vss 31.5253e-18
c849 n3__i5__i8__i10__net22 vss 76.9463e-18
c850 n3__i5__i6__i5__net22 vss 84.3487e-18
c851 n66__i1__net2 vss 14.3856e-18
c852 n68__i1__net2 vss 14.4137e-18
c853 n58__i1__net2 vss 44.2943e-18
c854 n60__i1__net2 vss 51.5398e-18
c855 n54__i1__net2 vss 60.5214e-18
c856 n56__i1__net2 vss 53.0435e-18
c857 n13__i5__i8__net1 vss 18.2615e-18
c858 n12__i5__i8__net2 vss 23.8755e-18
c859 n34__i5__i6__net31 vss 18.5805e-18
c860 n55__i5__clk_buf vss 24.6983e-18
c861 n50__i1__net2 vss 14.1998e-18
c862 n52__i1__net2 vss 14.228e-18
c863 n3__i5__i8__net5 vss 89.6595e-18
c864 n3__i5__i6__net35 vss 77.951e-18
c865 n46__i1__net2 vss 14.3856e-18
c866 n48__i1__net2 vss 14.4137e-18
c867 n42__i1__net2 vss 14.1998e-18
c868 n44__i1__net2 vss 14.228e-18
c869 n33__shift vss 204.503e-18
c870 n4__i5__i6__i8__net4 vss 221.269e-18
c871 n38__i1__net2 vss 14.3856e-18
c872 n40__i1__net2 vss 14.4137e-18
c873 n4__i5__i8__net2 vss 73.488e-18
c874 n34__i1__net2 vss 56.6537e-18
c875 n36__i1__net2 vss 52.9428e-18
c876 n2__i5__i6__i8__net4 vss 86.7068e-18
c877 n31__shift vss 229.119e-18
c878 n30__i1__net2 vss 60.8724e-18
c879 n32__i1__net2 vss 50.5187e-18
c880 n26__i1__net2 vss 14.1998e-18
c881 n28__i1__net2 vss 14.228e-18
c882 n24__shift vss 24.3469e-18
c883 n49__reset vss 31.6537e-18
c884 n22__i1__net2 vss 14.3856e-18
c885 n24__i1__net2 vss 14.4137e-18
c886 n18__i1__net2 vss 14.1247e-18
c887 n20__i1__net2 vss 14.1531e-18
c888 n7__i5__i8__net4 vss 208.389e-18
c889 n42__i5__clk_buf vss 26.9574e-18
c890 n14__i1__net2 vss 53.4922e-18
c891 n16__i1__net2 vss 62.8058e-18
c892 n45__reset vss 118.37e-18
c893 n3__i5__i8__i9__net22 vss 78.8789e-18
c894 n9__i1__net2 vss 14.1722e-18
c895 n11__i1__net2 vss 14.2004e-18
c896 n28__i5__i6__net31 vss 234.939e-18
c897 n39__i5__clk_buf vss 31.6559e-18
c898 n6__i1__net2 vss 14.5667e-18
c899 n8__i1__net2 vss 14.6097e-18
c900 n3__i5__i6__i4__net22 vss 80.252e-18
c901 n3__i1__net2 vss 21.6474e-18
c902 n3__i5__i8__net4 vss 18.1545e-18
c903 n34__i5__clk_buf vss 23.9803e-18
c904 n3__i5__i8__net1 vss 62.9237e-18
c905 n20__i5__i6__net31 vss 18.5805e-18
c906 n31__i5__clk_buf vss 25.8618e-18
c907 n3__i5__i6__net33 vss 76.3462e-18
c908 n21__i5__clk_buf vss 76.7622e-18
c909 n20__shift vss 202.801e-18
c910 n4__i5__i6__i7__net4 vss 220.826e-18
c911 n14__i5__i9__net21 vss 55.2265e-18
c912 n16__i5__i9__net21 vss 49.5153e-18
c913 n2__i5__i6__i7__net4 vss 87.9485e-18
c914 n18__shift vss 228.386e-18
c915 n10__i5__i9__net21 vss 71.4014e-18
c916 n12__i5__i9__net21 vss 56.9133e-18
c917 n6__i5__i9__net21 vss 62.8616e-18
c918 n8__i5__i9__net21 vss 57.3018e-18
c919 n714__i1__i14__net1 vss 22.4621e-18
c920 n716__i1__i14__net1 vss 21.9987e-18
c921 n5__i5__i9__net21 vss 51.8439e-18
c922 n3__i5__i9__net21 vss 118.081e-18
c923 n11__shift vss 23.4922e-18
c924 n706__i1__i14__net1 vss 14.5093e-18
c925 n708__i1__i14__net1 vss 14.3197e-18
c926 n702__i1__i14__net1 vss 14.2938e-18
c927 n704__i1__i14__net1 vss 14.1088e-18
c928 n4__clk_out vss 19.6445e-18
c929 n690__i1__i14__net1 vss 50.7988e-18
c930 n692__i1__i14__net1 vss 61.5362e-18
c931 n38__reset vss 32.9298e-18
c932 n686__i1__i14__net1 vss 60.9288e-18
c933 n688__i1__i14__net1 vss 49.9727e-18
c934 n2__i5__i7__i7__net3 vss 100.711e-18
c935 n674__i1__i14__net1 vss 14.4796e-18
c936 n676__i1__i14__net1 vss 14.9531e-18
c937 n7__i5__i6__net31 vss 236.064e-18
c938 n15__i5__clk_buf vss 31.6205e-18
c939 n670__i1__i14__net1 vss 14.2938e-18
c940 n672__i1__i14__net1 vss 14.1088e-18
c941 n3__i5__i6__i2__net22 vss 81.6147e-18
c942 n658__i1__i14__net1 vss 14.4045e-18
c943 n660__i1__i14__net1 vss 14.8783e-18
c944 n19__i5__i7__net44 vss 235.077e-18
c945 n17__i5__i7__i7__net1 vss 32.4926e-18
c946 n650__i1__i14__net1 vss 14.5935e-18
c947 n652__i1__i14__net1 vss 14.4056e-18
c948 n10__i5__i7__net46 vss 40.9083e-18
c949 n14__i5__i7__i7__net1 vss 155.098e-18
c950 n3__i5__i6__net31 vss 18.5805e-18
c951 n12__i5__clk_buf vss 102.067e-18
c952 n646__i1__i14__net1 vss 14.6814e-18
c953 n648__i1__i14__net1 vss 14.4901e-18
c954 n3__i5__i6__net30 vss 76.4658e-18
c955 n4__i5__i7__i7__net2 vss 155.265e-18
c956 n9__i5__i7__net46 vss 39.6807e-18
c957 n638__i1__i14__net1 vss 14.6814e-18
c958 n640__i1__i14__net1 vss 14.4901e-18
c959 n630__i1__i14__net1 vss 14.6814e-18
c960 n632__i1__i14__net1 vss 14.4901e-18
c961 n2__i5__i7__i7__net2 vss 30.4208e-18
c962 n11__i5__i7__net44 vss 33.6937e-18
c963 n7__shift vss 202.726e-18
c964 n4__i5__i6__i6__net4 vss 236.096e-18
c965 n618__i1__i14__net1 vss 14.6814e-18
c966 n620__i1__i14__net1 vss 14.4901e-18
c967 n610__i1__i14__net1 vss 14.6814e-18
c968 n612__i1__i14__net1 vss 15.1235e-18
c969 n2__i5__i6__i6__net4 vss 85.716e-18
c970 n5__shift vss 229.288e-18
c971 n606__i1__i14__net1 vss 14.6814e-18
c972 n608__i1__i14__net1 vss 14.4901e-18
c973 n7__i5__i7__i7__net1 vss 65.5221e-18
c974 n594__i1__i14__net1 vss 14.6814e-18
c975 n596__i1__i14__net1 vss 14.9613e-18
c976 n2__shift vss 25.1542e-18
c977 n590__i1__i14__net1 vss 53.9121e-18
c978 n592__i1__i14__net1 vss 62.1898e-18
c979 n5__i5__i7__i7__net1 vss 144.119e-18
c980 n2__i5__i7__i7__i1__net1 vss 161.897e-18
c981 n578__i1__i14__net1 vss 14.6814e-18
c982 n580__i1__i14__net1 vss 14.3395e-18
c983 n570__i1__i14__net1 vss 61.5015e-18
c984 n572__i1__i14__net1 vss 38.0138e-18
c985 n4__i5__clk_buf vss 60.9447e-18
c986 n2__i5__i7__net46 vss 168.332e-18
c987 n562__i1__i14__net1 vss 50.3988e-18
c988 n564__i1__i14__net1 vss 61.297e-18
c989 n554__i1__i14__net1 vss 61.5015e-18
c990 n556__i1__i14__net1 vss 37.0726e-18
c991 n7__i5__i7__net51 vss 157.1e-18
c992 n6__i5__i7__i6__net1 vss 33.3373e-18
c993 n546__i1__i14__net1 vss 14.6814e-18
c994 n548__i1__i14__net1 vss 14.3279e-18
c995 n2__i5__i7__i7__net1 vss 27.4633e-18
c996 n542__i1__i14__net1 vss 14.6541e-18
c997 n544__i1__i14__net1 vss 14.3163e-18
c998 n2__i5__i7__net50 vss 119.259e-18
c999 n530__i1__i14__net1 vss 50.1417e-18
c1000 n532__i1__i14__net1 vss 60.2162e-18
c1001 n4__i5__i7__net51 vss 140.842e-18
c1002 n526__i1__i14__net1 vss 14.3658e-18
c1003 n528__i1__i14__net1 vss 14.2448e-18
c1004 n5__i5__i7__net47 vss 154.097e-18
c1005 n2__i5__i7__i7__i0__net1 vss 169.085e-18
c1006 n514__i1__i14__net1 vss 14.2193e-18
c1007 n516__i1__i14__net1 vss 13.9582e-18
c1008 n3__i5__i7__i6__net1 vss 265.329e-18
c1009 n506__i1__i14__net1 vss 14.4796e-18
c1010 n508__i1__i14__net1 vss 14.9531e-18
c1011 n2__i5__i7__net44 vss 170.602e-18
c1012 n498__i1__i14__net1 vss 14.2938e-18
c1013 n500__i1__i14__net1 vss 13.9582e-18
c1014 n494__i1__i14__net1 vss 14.4796e-18
c1015 n496__i1__i14__net1 vss 15.5865e-18
c1016 n2__i5__i7__net47 vss 29.9886e-18
c1017 n2__i5__i7__net51 vss 28.0979e-18
c1018 n482__i1__i14__net1 vss 14.2938e-18
c1019 n484__i1__i14__net1 vss 13.9582e-18
c1020 n478__i1__i14__net1 vss 50.7988e-18
c1021 n480__i1__i14__net1 vss 60.7469e-18
c1022 n466__i1__i14__net1 vss 14.2938e-18
c1023 n468__i1__i14__net1 vss 13.9582e-18
c1024 n14__i5__i7__xor2 vss 155.466e-18
c1025 n6__i5__i7__i5__net1 vss 36.162e-18
c1026 n14__i5__i7__xor1 vss 157.558e-18
c1027 n6__i5__i7__i4__net1 vss 33.7536e-18
c1028 n458__i1__i14__net1 vss 14.4796e-18
c1029 n460__i1__i14__net1 vss 14.3197e-18
c1030 n450__i1__i14__net1 vss 14.2938e-18
c1031 n452__i1__i14__net1 vss 14.1088e-18
c1032 n2__i5__i7__xor3 vss 118.17e-18
c1033 n2__i5__i7__xor0 vss 117.676e-18
c1034 n442__i1__i14__net1 vss 14.4796e-18
c1035 n444__i1__i14__net1 vss 14.3197e-18
c1036 n434__i1__i14__net1 vss 14.2187e-18
c1037 n436__i1__i14__net1 vss 14.034e-18
c1038 n11__i5__i7__xor2 vss 145.609e-18
c1039 n11__i5__i7__xor1 vss 140.324e-18
c1040 n426__i1__i14__net1 vss 14.3917e-18
c1041 n428__i1__i14__net1 vss 14.8686e-18
c1042 n421__i1__i14__net1 vss 14.2663e-18
c1043 n423__i1__i14__net1 vss 14.1126e-18
c1044 n3__i5__i7__i5__net1 vss 42.9712e-18
c1045 n3__i5__i7__i4__net1 vss 42.9012e-18
c1046 n414__i1__i14__net1 vss 58.0796e-18
c1047 n416__i1__i14__net1 vss 51.9914e-18
c1048 n405__i1__i14__net1 vss 14.2663e-18
c1049 n407__i1__i14__net1 vss 14.1126e-18
c1050 n394__i1__i14__net1 vss 14.6548e-18
c1051 n396__i1__i14__net1 vss 14.5012e-18
c1052 n2__i5__i7__xor2 vss 29.0822e-18
c1053 n2__i5__i7__xor1 vss 28.9715e-18
c1054 n389__i1__i14__net1 vss 14.2663e-18
c1055 n391__i1__i14__net1 vss 14.1126e-18
c1056 n380__i1__i14__net1 vss 14.6548e-18
c1057 n382__i1__i14__net1 vss 14.5012e-18
c1058 n373__i1__i14__net1 vss 14.2663e-18
c1059 n375__i1__i14__net1 vss 14.1126e-18
c1060 n5__i5__i7__y3out vss 152.524e-18
c1061 n2__i5__i7__i9__net1 vss 157.756e-18
c1062 n12__i5__i7__y0out vss 150.766e-18
c1063 n2__i5__i7__i2__net1 vss 162.469e-18
c1064 n362__i1__i14__net1 vss 14.6548e-18
c1065 n364__i1__i14__net1 vss 14.5012e-18
c1066 n357__i1__i14__net1 vss 59.452e-18
c1067 n359__i1__i14__net1 vss 40.4794e-18
c1068 n2__i5__i7__x3out vss 171.89e-18
c1069 n9__i5__i7__x0out vss 172.282e-18
c1070 n346__i1__i14__net1 vss 15.2883e-18
c1071 n348__i1__i14__net1 vss 14.5012e-18
c1072 n341__i1__i14__net1 vss 14.2663e-18
c1073 n343__i1__i14__net1 vss 14.1126e-18
c1074 n2__i5__i7__y3out vss 28.2387e-18
c1075 n9__i5__i7__y0out vss 28.0567e-18
c1076 n334__i1__i14__net1 vss 58.38e-18
c1077 n336__i1__i14__net1 vss 54.4106e-18
c1078 n325__i1__i14__net1 vss 14.2663e-18
c1079 n327__i1__i14__net1 vss 14.1126e-18
c1080 n314__i1__i14__net1 vss 57.47e-18
c1081 n316__i1__i14__net1 vss 54.2678e-18
c1082 n12__i5__i7__y2out vss 148.008e-18
c1083 n2__i5__i7__i8__net1 vss 162.922e-18
c1084 n12__i5__i7__y1out vss 148.312e-18
c1085 n2__i5__i7__i3__net1 vss 165.881e-18
c1086 n305__i1__i14__net1 vss 14.3339e-18
c1087 n307__i1__i14__net1 vss 14.1799e-18
c1088 n302__i1__i14__net1 vss 15.3739e-18
c1089 n304__i1__i14__net1 vss 14.5834e-18
c1090 n2__i5__i7__x2out vss 170.744e-18
c1091 n9__i5__i7__x1out vss 171.034e-18
c1092 n294__i1__i14__net1 vss 14.2938e-18
c1093 n296__i1__i14__net1 vss 14.1088e-18
c1094 n286__i1__i14__net1 vss 50.9881e-18
c1095 n288__i1__i14__net1 vss 63.4349e-18
c1096 n2__i5__i7__y2out vss 27.7319e-18
c1097 n9__i5__i7__y1out vss 27.507e-18
c1098 n274__i1__i14__net1 vss 14.3729e-18
c1099 n276__i1__i14__net1 vss 14.1845e-18
c1100 n270__i1__i14__net1 vss 14.2047e-18
c1101 n272__i1__i14__net1 vss 14.5561e-18
c1102 n27__reset vss 62.5104e-18
c1103 n25__reset vss 60.6721e-18
c1104 n258__i1__i14__net1 vss 14.6814e-18
c1105 n260__i1__i14__net1 vss 14.4901e-18
c1106 n254__i1__i14__net1 vss 14.6814e-18
c1107 n256__i1__i14__net1 vss 14.4901e-18
c1108 n26__i5__i7__i1__net1 vss 79.3862e-18
c1109 n57__i5__clk4 vss 73.5166e-18
c1110 n26__i5__i7__i0__net1 vss 79.0625e-18
c1111 n55__i5__clk4 vss 69.0247e-18
c1112 n242__i1__i14__net1 vss 14.1384e-18
c1113 n244__i1__i14__net1 vss 14.4901e-18
c1114 n238__i1__i14__net1 vss 14.6814e-18
c1115 n240__i1__i14__net1 vss 14.4901e-18
c1116 n3__i5__i7__i1__i2__net22 vss 43.4877e-18
c1117 n3__i5__i7__i0__i2__net22 vss 43.2941e-18
c1118 n226__i1__i14__net1 vss 14.6814e-18
c1119 n228__i1__i14__net1 vss 14.4901e-18
c1120 n49__i5__clk4 vss 81.2101e-18
c1121 n22__i5__i7__i1__net1 vss 68.3683e-18
c1122 n47__i5__clk4 vss 83.1886e-18
c1123 n22__i5__i7__i0__net1 vss 67.006e-18
c1124 n218__i1__i14__net1 vss 14.6814e-18
c1125 n220__i1__i14__net1 vss 14.4901e-18
c1126 n210__i1__i14__net1 vss 14.0505e-18
c1127 n212__i1__i14__net1 vss 14.4056e-18
c1128 n3__y3 vss 7.86741e-18
c1129 n3__x3 vss 7.98077e-18
c1130 n202__i1__i14__net1 vss 53.4492e-18
c1131 n204__i1__i14__net1 vss 61.4775e-18
c1132 n198__i1__i14__net1 vss 14.2938e-18
c1133 n200__i1__i14__net1 vss 14.1088e-18
c1134 n19__reset vss 61.0977e-18
c1135 n17__reset vss 61.0328e-18
c1136 n186__i1__i14__net1 vss 53.5414e-18
c1137 n188__i1__i14__net1 vss 62.9588e-18
c1138 n178__i1__i14__net1 vss 14.2938e-18
c1139 n180__i1__i14__net1 vss 14.1088e-18
c1140 n19__i5__i7__i1__net1 vss 79.9849e-18
c1141 n43__i5__clk4 vss 73.2134e-18
c1142 n19__i5__i7__i0__net1 vss 82.5338e-18
c1143 n41__i5__clk4 vss 69.4647e-18
c1144 n174__i1__i14__net1 vss 14.4796e-18
c1145 n176__i1__i14__net1 vss 14.3197e-18
c1146 n3__i5__i7__i1__i1__net22 vss 42.4019e-18
c1147 n3__i5__i7__i0__i1__net22 vss 43.193e-18
c1148 n162__i1__i14__net1 vss 45.0051e-18
c1149 n164__i1__i14__net1 vss 52.808e-18
c1150 n158__i1__i14__net1 vss 14.4796e-18
c1151 n160__i1__i14__net1 vss 14.3197e-18
c1152 n39__i5__clk4 vss 81.1686e-18
c1153 n17__i5__i7__i1__net1 vss 67.7674e-18
c1154 n37__i5__clk4 vss 83.1744e-18
c1155 n17__i5__i7__i0__net1 vss 66.6272e-18
c1156 n146__i1__i14__net1 vss 14.2938e-18
c1157 n148__i1__i14__net1 vss 14.1088e-18
c1158 n142__i1__i14__net1 vss 53.5414e-18
c1159 n144__i1__i14__net1 vss 61.5699e-18
c1160 n3__y2 vss 8.02659e-18
c1161 n3__x2 vss 8.14083e-18
c1162 n132__i1__i14__net1 vss 14.2938e-18
c1163 n134__i1__i14__net1 vss 14.1088e-18
c1164 n8__reset vss 61.4722e-18
c1165 n6__reset vss 60.695e-18
c1166 n126__i1__i14__net1 vss 14.4796e-18
c1167 n128__i1__i14__net1 vss 14.3197e-18
c1168 n114__i1__i14__net1 vss 14.2938e-18
c1169 n116__i1__i14__net1 vss 14.1088e-18
c1170 n12__i5__i7__i1__net1 vss 78.8509e-18
c1171 n29__i5__clk4 vss 73.4447e-18
c1172 n12__i5__i7__i0__net1 vss 82.0239e-18
c1173 n27__i5__clk4 vss 69.8865e-18
c1174 n106__i1__i14__net1 vss 14.4796e-18
c1175 n108__i1__i14__net1 vss 14.3197e-18
c1176 n98__i1__i14__net1 vss 14.2938e-18
c1177 n100__i1__i14__net1 vss 14.1088e-18
c1178 n3__i5__i7__i1__i0__net22 vss 42.3393e-18
c1179 n3__i5__i7__i0__i0__net22 vss 42.3109e-18
c1180 n90__i1__i14__net1 vss 53.6717e-18
c1181 n92__i1__i14__net1 vss 59.2085e-18
c1182 n18__i5__clk4 vss 81.183e-18
c1183 n6__i5__i7__i1__net1 vss 68.1196e-18
c1184 n16__i5__clk4 vss 84.3424e-18
c1185 n6__i5__i7__i0__net1 vss 66.7792e-18
c1186 n82__i1__i14__net1 vss 43.5264e-18
c1187 n84__i1__i14__net1 vss 52.7517e-18
c1188 n78__i1__i14__net1 vss 14.3917e-18
c1189 n80__i1__i14__net1 vss 14.2352e-18
c1190 n3__y1 vss 8.19332e-18
c1191 n3__x1 vss 8.31459e-18
c1192 n65__i1__i14__net1 vss 14.2584e-18
c1193 n67__i1__i14__net1 vss 14.1126e-18
c1194 n58__i1__i14__net1 vss 53.6859e-18
c1195 n60__i1__i14__net1 vss 62.1718e-18
c1196 n4__reset vss 61.3236e-18
c1197 n2__reset vss 61.2132e-18
c1198 n53__i1__i14__net1 vss 14.1954e-18
c1199 n55__i1__i14__net1 vss 14.1126e-18
c1200 n50__i1__i14__net1 vss 14.585e-18
c1201 n52__i1__i14__net1 vss 14.5012e-18
c1202 n4__i5__i7__i1__net1 vss 81.1608e-18
c1203 n14__i5__clk4 vss 74.1249e-18
c1204 n4__i5__i7__i0__net1 vss 82.7654e-18
c1205 n12__i5__clk4 vss 70.2307e-18
c1206 n45__i1__i14__net1 vss 14.1954e-18
c1207 n47__i1__i14__net1 vss 14.1126e-18
c1208 n3__i5__i7__i1__i3__net22 vss 41.8819e-18
c1209 n3__i5__i7__i0__i3__net22 vss 42.0078e-18
c1210 n42__i1__i14__net1 vss 14.585e-18
c1211 n44__i1__i14__net1 vss 14.5012e-18
c1212 n37__i1__i14__net1 vss 14.1954e-18
c1213 n39__i1__i14__net1 vss 14.1126e-18
c1214 n10__i5__clk4 vss 80.5077e-18
c1215 n2__i5__i7__i1__net1 vss 68.32e-18
c1216 n8__i5__clk4 vss 82.4706e-18
c1217 n2__i5__i7__i0__net1 vss 66.9746e-18
c1218 n34__i1__i14__net1 vss 57.8158e-18
c1219 n36__i1__i14__net1 vss 54.0647e-18
c1220 n29__i1__i14__net1 vss 14.1954e-18
c1221 n31__i1__i14__net1 vss 14.1126e-18
c1222 n3__y0 vss 10.1924e-18
c1223 n3__x0 vss 10.3135e-18
c1224 n26__i1__i14__net1 vss 14.585e-18
c1225 n28__i1__i14__net1 vss 14.5012e-18
c1226 n21__i1__i14__net1 vss 14.119e-18
c1227 n23__i1__i14__net1 vss 14.0365e-18
c1228 n5__i5__clk4 vss 31.0104e-18
c1229 n2__i5__clk4 vss 26.0366e-18
c1230 n18__i1__i14__net1 vss 14.6855e-18
c1231 n20__i1__i14__net1 vss 14.5892e-18
c1232 n14__i1__i14__net1 vss 48.7333e-18
c1233 n16__i1__i14__net1 vss 41.1572e-18
c1234 n10__i1__i14__net1 vss 14.6341e-18
c1235 n12__i1__i14__net1 vss 14.5376e-18
c1236 n6__i1__i14__net1 vss 14.6976e-18
c1237 n8__i1__i14__net1 vss 15.0563e-18
c1238 n4__i1__i14__net1 vss 24.2718e-18
c1239 n2__i1__i14__net1 vss 24.2372e-18
c1240 n482__vdd vss 353.973e-18
c1241 n485__vdd vss 1.04211e-15
c1242 n2100__vddio vss 426.735e-18
c1243 n427__vdd vss 100.439e-18
c1244 n431__vdd vss 153.104e-18
c1245 n1720__vddio vss 14.4635e-18
c1246 n1722__vddio vss 233.642e-21
c1247 n421__vdd vss 107.968e-18
c1248 n425__vdd vss 194.998e-18
c1249 n1672__vddio vss 59.9715e-18
c1250 n1674__vddio vss 15.4208e-18
c1251 n1676__vddio vss 4.11981e-18
c1252 n175__vdd vss 116.411e-18
c1253 n179__vdd vss 188.908e-18
c1254 n1403__vddio vss 71.5628e-18
c1255 n1405__vddio vss 25.2829e-18
c1256 n1407__vddio vss 2.4817e-18
c1257 n169__vdd vss 111.579e-18
c1258 n173__vdd vss 176.638e-18
c1259 n1288__vddio vss 68.5704e-18
c1260 n1290__vddio vss 23.8417e-18
c1261 n1292__vddio vss 3.27238e-18
c1262 n163__vdd vss 121.068e-18
c1263 n167__vdd vss 204.785e-18
c1264 n1194__vddio vss 46.3139e-18
c1265 n1196__vddio vss 34.392e-18
c1266 n1198__vddio vss 4.94159e-18
c1267 n145__vdd vss 132.297e-18
c1268 n149__vdd vss 244.726e-18
c1269 n1026__vddio vss 36.4585e-18
c1270 n1028__vddio vss 2.7549e-18
c1271 n1030__vddio vss 4.54294e-18
c1272 n37__vdd vss 132.957e-18
c1273 n41__vdd vss 206.465e-18
c1274 n908__vddio vss 348.736e-18
c1275 n910__vddio vss 35.8052e-18
c1276 n912__vddio vss 304.191e-21
c1277 n1577__chipdriverout vss 614.515e-18
c1278 n31__vdd vss 135.893e-18
c1279 n35__vdd vss 199.211e-18
c1280 n821__vddio vss 189.717e-18
c1281 n823__vddio vss 5.02738e-18
c1282 n825__vddio vss 4.6076e-18
c1283 n25__vdd vss 131.928e-18
c1284 n29__vdd vss 193.877e-18
c1285 n643__vddio vss 71.4318e-18
c1286 n645__vddio vss 24.7436e-18
c1287 n647__vddio vss 4.52702e-18
c1288 n19__vdd vss 122.472e-18
c1289 n23__vdd vss 185.002e-18
c1290 n570__vddio vss 69.3421e-18
c1291 n572__vddio vss 24.376e-18
c1292 n574__vddio vss 341.519e-21
c1293 n13__vdd vss 122.821e-18
c1294 n17__vdd vss 207.061e-18
c1295 n459__vddio vss 4.56373e-18
c1296 n455__vddio vss 58.3474e-18
c1297 n7__vdd vss 131.052e-18
c1298 n11__vdd vss 201.277e-18
c1299 n277__vddio vss 70.79e-18
c1300 n279__vddio vss 24.6143e-18
c1301 n281__vddio vss 4.52537e-18
c1302 n3__vdd vss 228.363e-18
c1303 n89__vddio vss 6.14007e-18
c1304 n91__vddio vss 16.1608e-18
c1305 n93__vddio vss 1.8659e-18
c1306 n434__vdd vss 131.433e-18
c1307 n462__vdd vss 77.5256e-18
c1308 n478__vdd vss 201.823e-18
c1309 n2071__vddio vss 456.416e-21
c1310 n428__vdd vss 91.8145e-18
c1311 n429__vdd vss 66.22e-18
c1312 n432__vdd vss 203.678e-18
c1313 n422__vdd vss 67.4585e-18
c1314 n423__vdd vss 104.462e-18
c1315 n426__vdd vss 204.374e-18
c1316 n177__vdd vss 233.159e-18
c1317 n180__vdd vss 179.247e-18
c1318 n1408__vddio vss 9.04007e-21
c1319 n170__vdd vss 91.7439e-18
c1320 n171__vdd vss 244.548e-18
c1321 n174__vdd vss 280.118e-18
c1322 n164__vdd vss 45.3916e-18
c1323 n165__vdd vss 273.51e-18
c1324 n168__vdd vss 383.056e-18
c1325 n146__vdd vss 194.409e-18
c1326 n147__vdd vss 340.164e-18
c1327 n150__vdd vss 408.218e-18
c1328 n1031__vddio vss 9.83462e-21
c1329 n38__vdd vss 29.5534e-18
c1330 n39__vdd vss 257.647e-18
c1331 n42__vdd vss 309.008e-18
c1332 n913__vddio vss 9.04007e-21
c1333 n1537__chipdriverout vss 8.25471e-18
c1334 n32__vdd vss 28.8493e-18
c1335 n33__vdd vss 237.364e-18
c1336 n36__vdd vss 236.642e-18
c1337 n26__vdd vss 53.6282e-18
c1338 n27__vdd vss 223.676e-18
c1339 n30__vdd vss 235.638e-18
c1340 n20__vdd vss 33.1841e-18
c1341 n21__vdd vss 235.756e-18
c1342 n24__vdd vss 269.949e-18
c1343 n575__vddio vss 9.04007e-21
c1344 n14__vdd vss 39.5264e-18
c1345 n15__vdd vss 292.786e-18
c1346 n18__vdd vss 278.189e-18
c1347 n457__vddio vss 3.13376e-18
c1348 n460__vddio vss 8.24551e-21
c1349 n8__vdd vss 48.4109e-18
c1350 n9__vdd vss 315.416e-18
c1351 n12__vdd vss 296.521e-18
c1352 n282__vddio vss 14.1073e-21
c1353 n204__vddio vss 4.11604e-18
c1354 n206__vddio vss 25.298e-18
c1355 n208__vddio vss 50.1493e-21
c1356 n1__vdd vss 56.5795e-18
c1357 n5__vdd vss 206.453e-18
c1358 n94__vddio vss 1.58912e-21
c1359 n2024__vddio vss 12.4539e-18
c1360 n2023__vddio vss 16.1057e-18
c1361 n2020__vddio vss 13.771e-18
c1362 n2019__vddio vss 30.9912e-18
c1363 n1729__vddio vss 18.3202e-18
c1364 n1728__vddio vss 11.2793e-18
c1365 n1726__vddio vss 8.6473e-21
c1366 n1671__vddio vss 68.9626e-18
c1367 n1670__vddio vss 52.3733e-18
c1368 n1668__vddio vss 9.26314e-18
c1369 n412__vdd vss 37.258e-18
c1370 n1402__vddio vss 27.0176e-18
c1371 n1401__vddio vss 17.2168e-18
c1372 n1399__vddio vss 9.10468e-18
c1373 n416__vdd vss 15.0996e-18
c1374 n1284__vddio vss 28.6806e-18
c1375 n1285__vddio vss 18.5997e-18
c1376 n1286__vddio vss 9.4093e-18
c1377 n1172__vddio vss 99.2346e-18
c1378 n1171__vddio vss 78.5149e-18
c1379 n1169__vddio vss 7.30916e-18
c1380 n420__vdd vss 61.3332e-18
c1381 n1035__vddio vss 69.9343e-18
c1382 n1034__vddio vss 45.9133e-18
c1383 n1032__vddio vss 9.1505e-18
c1384 n125__vdd vss 37.4022e-18
c1385 n907__vddio vss 34.0984e-18
c1386 n906__vddio vss 24.3644e-18
c1387 n904__vddio vss 22.8003e-18
c1388 n1497__chipdriverout vss 997.991e-21
c1389 n796__vddio vss 125.507e-18
c1390 n797__vddio vss 47.9448e-18
c1391 n798__vddio vss 10.788e-21
c1392 n129__vdd vss 34.4181e-18
c1393 n642__vddio vss 28.452e-18
c1394 n641__vddio vss 18.2818e-18
c1395 n639__vddio vss 5.02398e-18
c1396 n566__vddio vss 27.7305e-18
c1397 n567__vddio vss 18.1367e-18
c1398 n425__vddio vss 52.6152e-18
c1399 n426__vddio vss 59.5947e-18
c1400 n137__vdd vss 32.825e-18
c1401 n276__vddio vss 28.2128e-18
c1402 n275__vddio vss 18.1314e-18
c1403 n273__vddio vss 3.81137e-18
c1404 n200__vddio vss 64.2139e-18
c1405 n201__vddio vss 17.7263e-18
c1406 n202__vddio vss 197.663e-21
c1407 n144__vdd vss 53.9008e-18
c1408 n64__vddio vss 47.7454e-18
c1409 n65__vddio vss 33.6063e-18
c1410 n66__vddio vss 725.945e-21
c1411 n1983__vddio vss 955.179e-24
c1412 n1986__vddio vss 955.179e-24
c1413 n403__vdd vss 12.4535e-18
c1414 n405__vdd vss 54.7568e-18
c1415 n17__i5__r0 vss 626.36e-18
c1416 n411__vdd vss 32.6533e-18
c1417 n15__i5__r1 vss 284.223e-18
c1418 n14__i5__r2 vss 355.552e-18
c1419 n9__i5__r1 vss 232.776e-18
c1420 n2__i5__r2 vss 261.345e-18
c1421 n3__i5__r0 vss 570.989e-18
c1422 n799__vddio vss 3.58708e-18
c1423 n110__vdd vss 13.8161e-18
c1424 n112__vdd vss 23.3583e-18
c1425 n568__vddio vss 22.4274e-18
c1426 n423__vddio vss 3.40634e-18
c1427 n118__vdd vss 24.7774e-18
c1428 n120__vdd vss 28.9761e-18
c1429 n122__vdd vss 28.244e-18
c1430 n203__vddio vss 22.3417e-18
c1431 n67__vddio vss 5.0528e-18
c1432 n1944__vddio vss 5.48505e-18
c1433 n1946__vddio vss 14.6798e-21
c1434 n1948__vddio vss 591.039e-18
c1435 n1950__vddio vss 6.33057e-18
c1436 n394__vdd vss 31.2245e-18
c1437 n1952__vddio vss 18.2356e-18
c1438 n40__i5__i8__net2 vss 246.241e-18
c1439 n396__vdd vss 55.9368e-18
c1440 n19__i5__i8__net2 vss 287.821e-18
c1441 n64__reset vss 221.889e-18
c1442 n67__reset vss 300.93e-18
c1443 n402__vdd vss 55.6401e-18
c1444 n14__i5__r1 vss 25.0426e-18
c1445 n13__i5__r2 vss 34.6001e-18
c1446 n8__i5__r1 vss 262.511e-18
c1447 n7__clk_out vss 239e-18
c1448 n1962__vddio vss 17.2728e-18
c1449 n2__i5__r0 vss 58.2947e-18
c1450 n1443__chipdriverout vss 127.434e-18
c1451 n1966__vddio vss 16.7285e-18
c1452 n90__vdd vss 33.4496e-18
c1453 n1970__vddio vss 14.7819e-18
c1454 n96__vdd vss 65.9696e-18
c1455 n98__vdd vss 52.1404e-18
c1456 n100__vdd vss 51.5746e-18
c1457 n1980__vddio vss 4.19839e-21
c1458 n13__reset vss 1.28836e-15
c1459 n105__vdd vss 23.4617e-18
c1460 n1982__vddio vss 18.14e-18
c1461 n21__i5__clk4 vss 2.02964e-15
c1462 n1892__vddio vss 24.1767e-18
c1463 n19__piso_outinv vss 450.375e-18
c1464 n1898__vddio vss 39.7545e-18
c1465 n30__piso_out vss 109.864e-18
c1466 n1904__vddio vss 33.4421e-18
c1467 n1737__vddio vss 1.70257e-15
c1468 n3__piso_outinv vss 451.944e-18
c1469 n39__i5__i8__net2 vss 3.94199e-18
c1470 n19__piso_out vss 434.364e-18
c1471 n99__i5__clk4 vss 2.24184e-15
c1472 n19__i5__i8__net5 vss 154.701e-18
c1473 n41__shift vss 966.579e-18
c1474 n72__reset vss 163.613e-18
c1475 n43__i5__i6__net31 vss 223.967e-18
c1476 n10__i5__i8__net5 vss 197.529e-18
c1477 n25__i5__i8__net1 vss 188.931e-18
c1478 n15__i5__r0 vss 13.0676e-18
c1479 n1915__vddio vss 4.19839e-21
c1480 n18__i5__i8__net2 vss 15.3863e-18
c1481 n37__shift vss 278.061e-18
c1482 n391__vdd vss 162.997e-18
c1483 n52__reset vss 298.091e-18
c1484 n10__i5__i8__net1 vss 209.802e-18
c1485 n31__i5__i6__net31 vss 28.673e-18
c1486 n778__i1__i14__net1 vss 128.061e-18
c1487 n779__i1__i14__net1 vss 104.342e-18
c1488 n780__i1__i14__net1 vss 115.392e-18
c1489 n781__i1__i14__net1 vss 104.617e-18
c1490 n782__i1__i14__net1 vss 103.808e-18
c1491 n783__i1__i14__net1 vss 65.5781e-18
c1492 n784__i1__i14__net1 vss 69.2223e-18
c1493 n785__i1__i14__net1 vss 71.3251e-18
c1494 n786__i1__i14__net1 vss 70.5408e-18
c1495 n787__i1__i14__net1 vss 71.4437e-18
c1496 n788__i1__i14__net1 vss 122.291e-18
c1497 n789__i1__i14__net1 vss 114.18e-18
c1498 n790__i1__i14__net1 vss 125.769e-18
c1499 n777__i1__i14__net1 vss 121.898e-18
c1500 n393__vdd vss 45.9276e-18
c1501 n13__i5__r1 vss 48.661e-18
c1502 n27__shift vss 29.1083e-18
c1503 n10__clk_out vss 130.103e-18
c1504 n42__reset vss 167.812e-18
c1505 n23__i5__i6__net31 vss 48.6291e-18
c1506 n67__vdd vss 110.58e-18
c1507 n14__shift vss 44.1031e-18
c1508 n16__i5__i6__net31 vss 226.089e-18
c1509 n7__i5__r1 vss 209.453e-18
c1510 n69__vdd vss 91.6079e-18
c1511 n1496__chipdriverout vss 291.691e-18
c1512 n1495__chipdriverout vss 296.116e-18
c1513 n1494__chipdriverout vss 325.223e-18
c1514 n1493__chipdriverout vss 300.06e-18
c1515 n1492__chipdriverout vss 188.41e-18
c1516 n1484__chipdriverout vss 198.968e-18
c1517 n1485__chipdriverout vss 238.762e-18
c1518 n1486__chipdriverout vss 277.074e-18
c1519 n1487__chipdriverout vss 242.257e-18
c1520 n1488__chipdriverout vss 250.872e-18
c1521 n1489__chipdriverout vss 296.884e-18
c1522 n1490__chipdriverout vss 316.996e-18
c1523 n1491__chipdriverout vss 258.592e-18
c1524 n71__vdd vss 55.0602e-18
c1525 n73__vdd vss 110.817e-18
c1526 n12__i5__i7__x3out vss 152.825e-18
c1527 n11__i5__i7__x0out vss 690.334e-18
c1528 n14__i5__i7__y0out vss 1.0848e-15
c1529 n77__vdd vss 55.6845e-18
c1530 n12__i5__i7__x2out vss 241.028e-18
c1531 n11__i5__i7__x1out vss 650.132e-18
c1532 n13__i5__i7__y2out vss 176.116e-18
c1533 n15__i5__i7__y1out vss 553.342e-18
c1534 n1933__vddio vss 5.43022e-21
c1535 n10__i5__i7__x3out vss 221.855e-18
c1536 n79__vdd vss 80.0718e-18
c1537 n10__i5__i7__y2out vss 241.324e-18
c1538 n10__i5__i7__x2out vss 202.129e-18
c1539 n81__vdd vss 82.1123e-18
c1540 n1937__vddio vss 5.43022e-21
c1541 n7__i5__i7__y1out vss 402.293e-18
c1542 n7__i5__i7__x1out vss 644.85e-18
c1543 n83__vdd vss 135.402e-18
c1544 n7__i5__i7__y0out vss 918.442e-18
c1545 n7__i5__i7__x0out vss 667.587e-18
c1546 n15__reset vss 253.749e-18
c1547 n14__reset vss 217.937e-18
c1548 n1941__vddio vss 3.52307e-21
c1549 n20__i5__clk4 vss 6.4693e-18
c1550 n78__i1__net3 vss 1.10502e-15
c1551 n1879__vddio vss 38.4955e-18
c1552 n76__i1__net3 vss 59.0401e-18
c1553 n74__i1__net3 vss 43.1909e-18
c1554 n72__i1__net3 vss 42.2003e-18
c1555 n70__i1__net3 vss 41.8504e-18
c1556 n66__i1__net3 vss 37.3183e-18
c1557 n67__i1__net3 vss 84.3696e-18
c1558 n209__i1__i13__net1 vss 193.399e-18
c1559 n212__i1__i13__net1 vss 218.334e-18
c1560 n202__i1__i13__net1 vss 195.547e-18
c1561 n205__i1__i13__net1 vss 151.214e-18
c1562 n206__i1__i13__net1 vss 212.932e-18
c1563 n200__i1__i13__net1 vss 13.8956e-18
c1564 n201__i1__i13__net1 vss 37.4497e-18
c1565 n18__piso_outinv vss 99.2016e-18
c1566 n1835__vddio vss 14.2987e-18
c1567 n196__i1__i13__net1 vss 16.9758e-18
c1568 n197__i1__i13__net1 vss 39.0798e-18
c1569 n192__i1__i13__net1 vss 39.276e-18
c1570 n193__i1__i13__net1 vss 39.0413e-18
c1571 n1883__vddio vss 22.7382e-18
c1572 n143__i1__i13__net1 vss 39.6548e-18
c1573 n144__i1__i13__net1 vss 38.2225e-18
c1574 n29__piso_out vss 61.2303e-18
c1575 n1841__vddio vss 5.32968e-18
c1576 n135__i1__i13__net1 vss 39.7828e-18
c1577 n136__i1__i13__net1 vss 39.6026e-18
c1578 n21__i1__net4 vss 93.7342e-18
c1579 n19__i1__net4 vss 51.506e-18
c1580 n127__i1__i13__net1 vss 43.2736e-18
c1581 n128__i1__i13__net1 vss 26.102e-18
c1582 n15__i1__net4 vss 105.522e-18
c1583 n115__i1__i13__net1 vss 71.8435e-18
c1584 n116__i1__i13__net1 vss 35.6204e-18
c1585 n1732__vddio vss 76.7513e-18
c1586 n57__i1__i12__net1 vss 146.288e-18
c1587 n1885__vddio vss 29.1073e-18
c1588 n105__i1__i13__net1 vss 39.3021e-18
c1589 n108__i1__i13__net1 vss 72.7544e-18
c1590 n51__i1__i12__net1 vss 66.9823e-18
c1591 n52__i1__i12__net1 vss 43.0454e-18
c1592 n93__i1__i13__net1 vss 63.3957e-18
c1593 n96__i1__i13__net1 vss 56.9135e-18
c1594 n44__i1__i12__net1 vss 51.7059e-18
c1595 n40__i1__i12__net1 vss 9.21729e-18
c1596 n75__i1__i13__net1 vss 39.258e-18
c1597 n76__i1__i13__net1 vss 87.6794e-18
c1598 n35__i1__i12__net1 vss 101.827e-18
c1599 n31__i1__i12__net1 vss 62.3785e-18
c1600 n32__i1__i12__net1 vss 24.4083e-18
c1601 n63__i1__i13__net1 vss 90.5139e-18
c1602 n64__i1__i13__net1 vss 43.2999e-18
c1603 n229__i1__net2 vss 248.853e-18
c1604 n228__i1__net2 vss 180.574e-18
c1605 n227__i1__net2 vss 202.422e-18
c1606 n226__i1__net2 vss 117.972e-18
c1607 n225__i1__net2 vss 114.518e-18
c1608 n1529__vddio vss 5.62749e-18
c1609 n1493__vddio vss 65.8098e-18
c1610 n1496__vddio vss 48.1706e-18
c1611 n1497__vddio vss 58.4879e-18
c1612 n1500__vddio vss 46.1649e-18
c1613 n1501__vddio vss 58.2357e-18
c1614 n1504__vddio vss 49.268e-18
c1615 n1505__vddio vss 52.65e-18
c1616 n1507__vddio vss 116.553e-18
c1617 n223__i1__net2 vss 281.93e-18
c1618 n1299__i1__i14__net1 vss 104.397e-18
c1619 n1300__i1__i14__net1 vss 85.386e-18
c1620 n1303__i1__i14__net1 vss 95.139e-18
c1621 n1304__i1__i14__net1 vss 82.5358e-18
c1622 n1307__i1__i14__net1 vss 55.9591e-18
c1623 n1308__i1__i14__net1 vss 105.002e-18
c1624 n1311__i1__i14__net1 vss 79.5867e-18
c1625 n1312__i1__i14__net1 vss 93.0647e-18
c1626 n1315__i1__i14__net1 vss 82.9441e-18
c1627 n1316__i1__i14__net1 vss 105.649e-18
c1628 n1319__i1__i14__net1 vss 90.7266e-18
c1629 n1320__i1__i14__net1 vss 118.556e-18
c1630 n1323__i1__i14__net1 vss 89.3903e-18
c1631 n219__i1__net2 vss 37.1748e-18
c1632 n1472__vddio vss 121.001e-18
c1633 n1475__vddio vss 119.256e-18
c1634 n1476__vddio vss 120.002e-18
c1635 n1479__vddio vss 121.524e-18
c1636 n1480__vddio vss 120.204e-18
c1637 n1483__vddio vss 114.381e-18
c1638 n1484__vddio vss 116.223e-18
c1639 n1508__vddio vss 77.7684e-18
c1640 n213__i1__net2 vss 37.6739e-18
c1641 n1285__i1__i14__net1 vss 117.448e-18
c1642 n1286__i1__i14__net1 vss 124.494e-18
c1643 n1287__i1__i14__net1 vss 136.635e-18
c1644 n1288__i1__i14__net1 vss 124.793e-18
c1645 n1289__i1__i14__net1 vss 93.3329e-18
c1646 n1290__i1__i14__net1 vss 91.3885e-18
c1647 n1291__i1__i14__net1 vss 119.849e-18
c1648 n1292__i1__i14__net1 vss 135.288e-18
c1649 n1293__i1__i14__net1 vss 120.055e-18
c1650 n1294__i1__i14__net1 vss 105.266e-18
c1651 n1295__i1__i14__net1 vss 125.884e-18
c1652 n1296__i1__i14__net1 vss 120.452e-18
c1653 n1297__i1__i14__net1 vss 127.855e-18
c1654 n38__i5__i8__net2 vss 35.9213e-18
c1655 n211__i1__net2 vss 37.3908e-18
c1656 n18__piso_out vss 15.8974e-18
c1657 n1465__vddio vss 103.698e-18
c1658 n1466__vddio vss 135.654e-18
c1659 n1467__vddio vss 104.319e-18
c1660 n1468__vddio vss 105.604e-18
c1661 n1469__vddio vss 104.319e-18
c1662 n1470__vddio vss 130.728e-18
c1663 n1471__vddio vss 100.526e-18
c1664 n1509__vddio vss 54.3615e-18
c1665 n207__i1__net2 vss 38.2475e-18
c1666 n98__i5__clk4 vss 78.0032e-18
c1667 n1246__i1__i14__net1 vss 126.511e-18
c1668 n1247__i1__i14__net1 vss 125.449e-18
c1669 n1248__i1__i14__net1 vss 137.288e-18
c1670 n1249__i1__i14__net1 vss 125.584e-18
c1671 n1250__i1__i14__net1 vss 92.9015e-18
c1672 n1251__i1__i14__net1 vss 91.557e-18
c1673 n1252__i1__i14__net1 vss 120.215e-18
c1674 n1253__i1__i14__net1 vss 135.621e-18
c1675 n1254__i1__i14__net1 vss 120.423e-18
c1676 n1255__i1__i14__net1 vss 105.698e-18
c1677 n1256__i1__i14__net1 vss 126.271e-18
c1678 n1257__i1__i14__net1 vss 120.875e-18
c1679 n1258__i1__i14__net1 vss 127.94e-18
c1680 n12__i5__i8__net5 vss 13.2758e-18
c1681 n203__i1__net2 vss 36.68e-18
c1682 n1444__vddio vss 121.584e-18
c1683 n1445__vddio vss 119.431e-18
c1684 n1446__vddio vss 120.406e-18
c1685 n1447__vddio vss 121.934e-18
c1686 n1448__vddio vss 120.609e-18
c1687 n1449__vddio vss 114.504e-18
c1688 n1450__vddio vss 116.597e-18
c1689 n1510__vddio vss 77.8356e-18
c1690 n199__i1__net2 vss 37.2803e-18
c1691 n1207__i1__i14__net1 vss 120.317e-18
c1692 n1208__i1__i14__net1 vss 108.877e-18
c1693 n1209__i1__i14__net1 vss 120.85e-18
c1694 n1210__i1__i14__net1 vss 107.392e-18
c1695 n1211__i1__i14__net1 vss 73.5267e-18
c1696 n1212__i1__i14__net1 vss 113.996e-18
c1697 n1213__i1__i14__net1 vss 104.506e-18
c1698 n1214__i1__i14__net1 vss 119.557e-18
c1699 n1215__i1__i14__net1 vss 104.506e-18
c1700 n1216__i1__i14__net1 vss 121.785e-18
c1701 n1217__i1__i14__net1 vss 111.512e-18
c1702 n1218__i1__i14__net1 vss 137.248e-18
c1703 n1219__i1__i14__net1 vss 111.898e-18
c1704 n40__shift vss 218.503e-18
c1705 n195__i1__net2 vss 43.79e-18
c1706 n378__vdd vss 172.339e-18
c1707 n1423__vddio vss 103.585e-18
c1708 n1424__vddio vss 135.669e-18
c1709 n1425__vddio vss 104.322e-18
c1710 n1426__vddio vss 105.603e-18
c1711 n1427__vddio vss 104.322e-18
c1712 n1428__vddio vss 130.796e-18
c1713 n1429__vddio vss 100.559e-18
c1714 n1511__vddio vss 54.6587e-18
c1715 n191__i1__net2 vss 36.8266e-18
c1716 n1168__i1__i14__net1 vss 103.873e-18
c1717 n1169__i1__i14__net1 vss 124.829e-18
c1718 n1170__i1__i14__net1 vss 137.103e-18
c1719 n1171__i1__i14__net1 vss 123.408e-18
c1720 n1172__i1__i14__net1 vss 90.6611e-18
c1721 n1173__i1__i14__net1 vss 90.9826e-18
c1722 n1174__i1__i14__net1 vss 119.893e-18
c1723 n1175__i1__i14__net1 vss 135.416e-18
c1724 n1176__i1__i14__net1 vss 120.098e-18
c1725 n1177__i1__i14__net1 vss 106.383e-18
c1726 n1178__i1__i14__net1 vss 130.459e-18
c1727 n1179__i1__i14__net1 vss 125.009e-18
c1728 n1180__i1__i14__net1 vss 126.045e-18
c1729 n186__i1__net2 vss 34.1931e-18
c1730 n1392__vddio vss 103.469e-18
c1731 n1393__vddio vss 135.525e-18
c1732 n1394__vddio vss 120.002e-18
c1733 n1395__vddio vss 121.524e-18
c1734 n1396__vddio vss 104.167e-18
c1735 n1397__vddio vss 129.154e-18
c1736 n1398__vddio vss 97.6638e-18
c1737 n1512__vddio vss 75.6793e-18
c1738 n71__reset vss 254.641e-18
c1739 n70__reset vss 14.2857e-18
c1740 n179__i1__net2 vss 35.1958e-18
c1741 n1129__i1__i14__net1 vss 120.11e-18
c1742 n1130__i1__i14__net1 vss 108.964e-18
c1743 n1131__i1__i14__net1 vss 120.849e-18
c1744 n1132__i1__i14__net1 vss 107.365e-18
c1745 n1133__i1__i14__net1 vss 72.5401e-18
c1746 n1134__i1__i14__net1 vss 114.355e-18
c1747 n1135__i1__i14__net1 vss 103.979e-18
c1748 n1136__i1__i14__net1 vss 118.98e-18
c1749 n1137__i1__i14__net1 vss 103.979e-18
c1750 n1138__i1__i14__net1 vss 124.939e-18
c1751 n1139__i1__i14__net1 vss 113.892e-18
c1752 n1140__i1__i14__net1 vss 139.133e-18
c1753 n1141__i1__i14__net1 vss 107.404e-18
c1754 n175__i1__net2 vss 34.4899e-18
c1755 n36__i5__i8__net2 vss 138.143e-18
c1756 n68__i5__clk_buf vss 105.002e-18
c1757 n1538__vddio vss 5.41914e-18
c1758 n1371__vddio vss 121.445e-18
c1759 n1372__vddio vss 119.248e-18
c1760 n1373__vddio vss 120.292e-18
c1761 n1374__vddio vss 121.819e-18
c1762 n1375__vddio vss 120.494e-18
c1763 n1376__vddio vss 113.727e-18
c1764 n1377__vddio vss 114.851e-18
c1765 n1513__vddio vss 77.0775e-18
c1766 n173__i1__net2 vss 36.8798e-18
c1767 n1065__i1__i14__net1 vss 120.449e-18
c1768 n1066__i1__i14__net1 vss 108.971e-18
c1769 n1069__i1__i14__net1 vss 120.85e-18
c1770 n1070__i1__i14__net1 vss 107.36e-18
c1771 n1073__i1__i14__net1 vss 72.9464e-18
c1772 n1074__i1__i14__net1 vss 114.247e-18
c1773 n1077__i1__i14__net1 vss 104.407e-18
c1774 n1078__i1__i14__net1 vss 119.374e-18
c1775 n1081__i1__i14__net1 vss 104.408e-18
c1776 n1082__i1__i14__net1 vss 121.748e-18
c1777 n1085__i1__i14__net1 vss 112.553e-18
c1778 n1086__i1__i14__net1 vss 139.124e-18
c1779 n1089__i1__i14__net1 vss 111.862e-18
c1780 n165__i1__net2 vss 37.4815e-18
c1781 n1337__vddio vss 101.845e-18
c1782 n1338__vddio vss 133.55e-18
c1783 n1341__vddio vss 102.49e-18
c1784 n1342__vddio vss 103.757e-18
c1785 n1345__vddio vss 102.49e-18
c1786 n1346__vddio vss 128.71e-18
c1787 n1349__vddio vss 98.7469e-18
c1788 n1514__vddio vss 53.6139e-18
c1789 n161__i1__net2 vss 36.9065e-18
c1790 n42__i5__i6__net31 vss 39.1454e-18
c1791 n1051__i1__i14__net1 vss 139.423e-18
c1792 n1052__i1__i14__net1 vss 108.51e-18
c1793 n1053__i1__i14__net1 vss 135.162e-18
c1794 n1054__i1__i14__net1 vss 108.328e-18
c1795 n1055__i1__i14__net1 vss 73.2918e-18
c1796 n1056__i1__i14__net1 vss 112.108e-18
c1797 n1057__i1__i14__net1 vss 102.596e-18
c1798 n1058__i1__i14__net1 vss 117.511e-18
c1799 n1059__i1__i14__net1 vss 102.596e-18
c1800 n1060__i1__i14__net1 vss 119.846e-18
c1801 n1061__i1__i14__net1 vss 108.561e-18
c1802 n1062__i1__i14__net1 vss 135.184e-18
c1803 n1063__i1__i14__net1 vss 109.811e-18
c1804 n66__i5__clk_buf vss 303.149e-18
c1805 n159__i1__net2 vss 40.3182e-18
c1806 n9__i5__i8__net5 vss 76.2787e-18
c1807 n1329__vddio vss 119.657e-18
c1808 n1330__vddio vss 117.847e-18
c1809 n1331__vddio vss 118.593e-18
c1810 n1332__vddio vss 120.096e-18
c1811 n1333__vddio vss 118.796e-18
c1812 n1334__vddio vss 113.011e-18
c1813 n1335__vddio vss 114.837e-18
c1814 n1515__vddio vss 53.7754e-18
c1815 n151__i1__net2 vss 41.1376e-18
c1816 n1012__i1__i14__net1 vss 140.361e-18
c1817 n1013__i1__i14__net1 vss 108.928e-18
c1818 n1014__i1__i14__net1 vss 119.482e-18
c1819 n1015__i1__i14__net1 vss 108.859e-18
c1820 n1016__i1__i14__net1 vss 73.3197e-18
c1821 n1017__i1__i14__net1 vss 112.607e-18
c1822 n1018__i1__i14__net1 vss 102.054e-18
c1823 n1019__i1__i14__net1 vss 116.804e-18
c1824 n1020__i1__i14__net1 vss 102.054e-18
c1825 n1021__i1__i14__net1 vss 119.553e-18
c1826 n1022__i1__i14__net1 vss 107.997e-18
c1827 n1023__i1__i14__net1 vss 134.684e-18
c1828 n1024__i1__i14__net1 vss 109.353e-18
c1829 n24__i5__i8__net1 vss 16.0413e-18
c1830 n143__i1__net2 vss 35.0984e-18
c1831 n1308__vddio vss 103.453e-18
c1832 n1309__vddio vss 135.503e-18
c1833 n1310__vddio vss 104.188e-18
c1834 n1311__vddio vss 105.471e-18
c1835 n1312__vddio vss 104.188e-18
c1836 n1313__vddio vss 130.628e-18
c1837 n1314__vddio vss 100.268e-18
c1838 n1516__vddio vss 76.8588e-18
c1839 n14__i5__r0 vss 18.8158e-18
c1840 n131__i1__net2 vss 35.7911e-18
c1841 n973__i1__i14__net1 vss 120.417e-18
c1842 n974__i1__i14__net1 vss 109.543e-18
c1843 n975__i1__i14__net1 vss 121.112e-18
c1844 n976__i1__i14__net1 vss 107.904e-18
c1845 n977__i1__i14__net1 vss 72.4499e-18
c1846 n978__i1__i14__net1 vss 114.047e-18
c1847 n979__i1__i14__net1 vss 104.13e-18
c1848 n980__i1__i14__net1 vss 119.168e-18
c1849 n981__i1__i14__net1 vss 104.13e-18
c1850 n982__i1__i14__net1 vss 123.03e-18
c1851 n983__i1__i14__net1 vss 115.14e-18
c1852 n984__i1__i14__net1 vss 141.698e-18
c1853 n985__i1__i14__net1 vss 109.438e-18
c1854 n125__i1__net2 vss 36.4599e-18
c1855 n1543__vddio vss 5.29959e-18
c1856 n1277__vddio vss 121.111e-18
c1857 n1278__vddio vss 119.418e-18
c1858 n1279__vddio vss 120.138e-18
c1859 n1280__vddio vss 121.661e-18
c1860 n1281__vddio vss 120.339e-18
c1861 n1282__vddio vss 113.241e-18
c1862 n1283__vddio vss 112.68e-18
c1863 n1517__vddio vss 75.9439e-18
c1864 n16__i5__i8__net2 vss 43.5506e-18
c1865 n117__i1__net2 vss 38.0394e-18
c1866 n934__i1__i14__net1 vss 120.343e-18
c1867 n935__i1__i14__net1 vss 109.536e-18
c1868 n936__i1__i14__net1 vss 121.112e-18
c1869 n937__i1__i14__net1 vss 107.908e-18
c1870 n938__i1__i14__net1 vss 72.4433e-18
c1871 n939__i1__i14__net1 vss 114.257e-18
c1872 n940__i1__i14__net1 vss 104.489e-18
c1873 n941__i1__i14__net1 vss 119.505e-18
c1874 n942__i1__i14__net1 vss 104.489e-18
c1875 n943__i1__i14__net1 vss 125.032e-18
c1876 n944__i1__i14__net1 vss 115.47e-18
c1877 n945__i1__i14__net1 vss 142.002e-18
c1878 n946__i1__i14__net1 vss 108.964e-18
c1879 n111__i1__net2 vss 34.1942e-18
c1880 n36__shift vss 99.2373e-18
c1881 n1242__vddio vss 121.493e-18
c1882 n1245__vddio vss 119.383e-18
c1883 n1246__vddio vss 120.349e-18
c1884 n1249__vddio vss 121.875e-18
c1885 n1250__vddio vss 120.551e-18
c1886 n1253__vddio vss 114.024e-18
c1887 n1254__vddio vss 115.221e-18
c1888 n1518__vddio vss 76.9038e-18
c1889 n55__reset vss 235.358e-18
c1890 n99__i1__net2 vss 45.4702e-18
c1891 n895__i1__i14__net1 vss 120.632e-18
c1892 n896__i1__i14__net1 vss 125.536e-18
c1893 n897__i1__i14__net1 vss 121.112e-18
c1894 n898__i1__i14__net1 vss 124.111e-18
c1895 n899__i1__i14__net1 vss 92.246e-18
c1896 n900__i1__i14__net1 vss 91.472e-18
c1897 n901__i1__i14__net1 vss 120.42e-18
c1898 n902__i1__i14__net1 vss 135.798e-18
c1899 n903__i1__i14__net1 vss 120.638e-18
c1900 n904__i1__i14__net1 vss 105.685e-18
c1901 n905__i1__i14__net1 vss 127.425e-18
c1902 n906__i1__i14__net1 vss 120.823e-18
c1903 n907__i1__i14__net1 vss 128.393e-18
c1904 n91__i1__net2 vss 35.8267e-18
c1905 n382__vdd vss 110.709e-18
c1906 n1235__vddio vss 103.625e-18
c1907 n1236__vddio vss 135.606e-18
c1908 n1237__vddio vss 104.261e-18
c1909 n1238__vddio vss 105.545e-18
c1910 n1239__vddio vss 104.261e-18
c1911 n1240__vddio vss 130.678e-18
c1912 n1241__vddio vss 100.467e-18
c1913 n1519__vddio vss 77.3463e-18
c1914 n64__i5__clk_buf vss 89.6519e-18
c1915 n82__i1__net2 vss 35.9871e-18
c1916 n51__reset vss 15.5054e-18
c1917 n856__i1__i14__net1 vss 142.198e-18
c1918 n857__i1__i14__net1 vss 110.707e-18
c1919 n858__i1__i14__net1 vss 121.703e-18
c1920 n859__i1__i14__net1 vss 110.643e-18
c1921 n860__i1__i14__net1 vss 74.108e-18
c1922 n861__i1__i14__net1 vss 114.333e-18
c1923 n862__i1__i14__net1 vss 104.038e-18
c1924 n863__i1__i14__net1 vss 118.992e-18
c1925 n864__i1__i14__net1 vss 104.038e-18
c1926 n865__i1__i14__net1 vss 121.616e-18
c1927 n866__i1__i14__net1 vss 110.068e-18
c1928 n867__i1__i14__net1 vss 136.947e-18
c1929 n868__i1__i14__net1 vss 111.601e-18
c1930 n79__i1__net2 vss 35.0629e-18
c1931 n1214__vddio vss 121.003e-18
c1932 n1215__vddio vss 119.234e-18
c1933 n1216__vddio vss 120.023e-18
c1934 n1217__vddio vss 121.547e-18
c1935 n1218__vddio vss 120.225e-18
c1936 n1219__vddio vss 114.361e-18
c1937 n1220__vddio vss 116.245e-18
c1938 n1520__vddio vss 54.2625e-18
c1939 n59__i5__clk_buf vss 96.619e-18
c1940 n71__i1__net2 vss 48.6251e-18
c1941 n817__i1__i14__net1 vss 160.125e-18
c1942 n818__i1__i14__net1 vss 139.477e-18
c1943 n819__i1__i14__net1 vss 157.808e-18
c1944 n820__i1__i14__net1 vss 140.488e-18
c1945 n821__i1__i14__net1 vss 94.7505e-18
c1946 n822__i1__i14__net1 vss 140.699e-18
c1947 n823__i1__i14__net1 vss 135.321e-18
c1948 n824__i1__i14__net1 vss 154.011e-18
c1949 n825__i1__i14__net1 vss 135.292e-18
c1950 n826__i1__i14__net1 vss 157.234e-18
c1951 n827__i1__i14__net1 vss 143.099e-18
c1952 n828__i1__i14__net1 vss 176.407e-18
c1953 n829__i1__i14__net1 vss 144.76e-18
c1954 n63__i1__net2 vss 55.4114e-18
c1955 n57__i5__clk_buf vss 212.118e-18
c1956 n1187__vddio vss 109.525e-18
c1957 n1188__vddio vss 100.92e-18
c1958 n1189__vddio vss 109.143e-18
c1959 n1190__vddio vss 110.362e-18
c1960 n1191__vddio vss 109.344e-18
c1961 n1192__vddio vss 95.2278e-18
c1962 n1193__vddio vss 105.042e-18
c1963 n8__i5__i8__net1 vss 55.337e-18
c1964 n30__i5__i6__net31 vss 40.5668e-18
c1965 n52__i5__clk_buf vss 49.9164e-18
c1966 n43__i5__clk_buf vss 147.981e-18
c1967 n1113__vddio vss 40.942e-18
c1968 n1114__vddio vss 28.6297e-18
c1969 n1115__vddio vss 30.1238e-18
c1970 n1116__vddio vss 30.4402e-18
c1971 n1117__vddio vss 29.7914e-18
c1972 n1118__vddio vss 32.8108e-18
c1973 n1119__vddio vss 30.8373e-18
c1974 n775__i1__i14__net1 vss 88.1198e-18
c1975 n1916__chipdriverout vss 104.039e-18
c1976 n1917__chipdriverout vss 83.7102e-18
c1977 n1918__chipdriverout vss 94.7881e-18
c1978 n1919__chipdriverout vss 83.4925e-18
c1979 n1920__chipdriverout vss 61.8523e-18
c1980 n1921__chipdriverout vss 96.7629e-18
c1981 n1922__chipdriverout vss 75.6138e-18
c1982 n1923__chipdriverout vss 85.8642e-18
c1983 n1924__chipdriverout vss 75.6139e-18
c1984 n1925__chipdriverout vss 97.4277e-18
c1985 n1926__chipdriverout vss 82.7636e-18
c1986 n1927__chipdriverout vss 112.081e-18
c1987 n1928__chipdriverout vss 87.5924e-18
c1988 n26__shift vss 97.0447e-18
c1989 n1551__vddio vss 6.77184e-18
c1990 n771__i1__i14__net1 vss 38.7495e-18
c1991 n1092__vddio vss 119.548e-18
c1992 n1093__vddio vss 117.243e-18
c1993 n1094__vddio vss 118.363e-18
c1994 n1095__vddio vss 119.871e-18
c1995 n1096__vddio vss 118.566e-18
c1996 n1097__vddio vss 112.406e-18
c1997 n1098__vddio vss 114.606e-18
c1998 n1121__vddio vss 77.3614e-18
c1999 n767__i1__i14__net1 vss 39.2646e-18
c2000 n1877__chipdriverout vss 141.292e-18
c2001 n1878__chipdriverout vss 109.885e-18
c2002 n1879__chipdriverout vss 121.526e-18
c2003 n1880__chipdriverout vss 109.126e-18
c2004 n1881__chipdriverout vss 76.4397e-18
c2005 n1882__chipdriverout vss 113.012e-18
c2006 n1883__chipdriverout vss 102.305e-18
c2007 n1884__chipdriverout vss 117.194e-18
c2008 n1885__chipdriverout vss 102.305e-18
c2009 n1886__chipdriverout vss 119.651e-18
c2010 n1887__chipdriverout vss 108.268e-18
c2011 n1888__chipdriverout vss 134.96e-18
c2012 n1889__chipdriverout vss 109.446e-18
c2013 n9__clk_out vss 28.4948e-18
c2014 n762__i1__i14__net1 vss 36.029e-18
c2015 n1071__vddio vss 102.383e-18
c2016 n1072__vddio vss 134.491e-18
c2017 n1073__vddio vss 103.174e-18
c2018 n1074__vddio vss 104.443e-18
c2019 n1075__vddio vss 103.174e-18
c2020 n1076__vddio vss 129.657e-18
c2021 n1077__vddio vss 99.8013e-18
c2022 n1122__vddio vss 54.3695e-18
c2023 n41__reset vss 24.4431e-18
c2024 n757__i1__i14__net1 vss 29.2469e-18
c2025 n8__i5__r2 vss 50.4974e-18
c2026 n1843__chipdriverout vss 90.9737e-18
c2027 n1844__chipdriverout vss 102.606e-18
c2028 n1845__chipdriverout vss 117.498e-18
c2029 n1846__chipdriverout vss 102.606e-18
c2030 n1847__chipdriverout vss 103.889e-18
c2031 n1848__chipdriverout vss 125.378e-18
c2032 n1849__chipdriverout vss 119.016e-18
c2033 n1850__chipdriverout vss 110.659e-18
c2034 n1813__chipdriverout vss 118.657e-18
c2035 n1814__chipdriverout vss 122.546e-18
c2036 n1817__chipdriverout vss 119.52e-18
c2037 n1818__chipdriverout vss 105.37e-18
c2038 n1821__chipdriverout vss 74.2627e-18
c2039 n755__i1__i14__net1 vss 36.9545e-18
c2040 n1050__vddio vss 105.615e-18
c2041 n1051__vddio vss 137.734e-18
c2042 n1052__vddio vss 106.181e-18
c2043 n1053__vddio vss 107.488e-18
c2044 n1054__vddio vss 106.181e-18
c2045 n1055__vddio vss 132.771e-18
c2046 n1056__vddio vss 102.05e-18
c2047 n1123__vddio vss 78.104e-18
c2048 n36__i5__clk_buf vss 96.0967e-18
c2049 n751__i1__i14__net1 vss 36.7757e-18
c2050 n1799__chipdriverout vss 103.453e-18
c2051 n1800__chipdriverout vss 123.889e-18
c2052 n1801__chipdriverout vss 137.09e-18
c2053 n1802__chipdriverout vss 122.705e-18
c2054 n1803__chipdriverout vss 92.1965e-18
c2055 n1804__chipdriverout vss 93.836e-18
c2056 n1805__chipdriverout vss 121.928e-18
c2057 n1806__chipdriverout vss 137.524e-18
c2058 n1807__chipdriverout vss 122.136e-18
c2059 n1808__chipdriverout vss 109.301e-18
c2060 n1809__chipdriverout vss 132.759e-18
c2061 n1810__chipdriverout vss 127.873e-18
c2062 n1811__chipdriverout vss 127.787e-18
c2063 n747__i1__i14__net1 vss 34.8456e-18
c2064 n1006__vddio vss 104.571e-18
c2065 n1007__vddio vss 136.594e-18
c2066 n1010__vddio vss 105.17e-18
c2067 n1011__vddio vss 106.465e-18
c2068 n1014__vddio vss 105.17e-18
c2069 n1015__vddio vss 129.696e-18
c2070 n1018__vddio vss 97.9257e-18
c2071 n1124__vddio vss 54.7478e-18
c2072 n28__i5__i7__i7__net1 vss 126.849e-18
c2073 n743__i1__i14__net1 vss 28.2957e-18
c2074 n1760__chipdriverout vss 120.714e-18
c2075 n1761__chipdriverout vss 108.634e-18
c2076 n1762__chipdriverout vss 121.649e-18
c2077 n1763__chipdriverout vss 107.221e-18
c2078 n1764__chipdriverout vss 74.256e-18
c2079 n1765__chipdriverout vss 115.693e-18
c2080 n1766__chipdriverout vss 105.089e-18
c2081 n1767__chipdriverout vss 120.158e-18
c2082 n1768__chipdriverout vss 105.09e-18
c2083 n1769__chipdriverout vss 125.269e-18
c2084 n1770__chipdriverout vss 116.179e-18
c2085 n1771__chipdriverout vss 142.522e-18
c2086 n1772__chipdriverout vss 109.863e-18
c2087 n22__i5__i6__net31 vss 16.4605e-18
c2088 n27__i5__clk_buf vss 274.306e-18
c2089 n739__i1__i14__net1 vss 37.7292e-18
c2090 n998__vddio vss 102.748e-18
c2091 n999__vddio vss 134.564e-18
c2092 n1000__vddio vss 103.372e-18
c2093 n1001__vddio vss 104.648e-18
c2094 n1002__vddio vss 103.372e-18
c2095 n1003__vddio vss 129.432e-18
c2096 n1004__vddio vss 98.5569e-18
c2097 n1125__vddio vss 53.8655e-18
c2098 n735__i1__i14__net1 vss 37.5438e-18
c2099 n19__i5__i7__net46 vss 221.786e-18
c2100 n1721__chipdriverout vss 102.275e-18
c2101 n1722__chipdriverout vss 122.561e-18
c2102 n1723__chipdriverout vss 136.042e-18
c2103 n1724__chipdriverout vss 121.549e-18
c2104 n1725__chipdriverout vss 92.8881e-18
c2105 n1726__chipdriverout vss 91.3182e-18
c2106 n1727__chipdriverout vss 119.006e-18
c2107 n1728__chipdriverout vss 134.332e-18
c2108 n1729__chipdriverout vss 119.213e-18
c2109 n1730__chipdriverout vss 104.416e-18
c2110 n1731__chipdriverout vss 125.963e-18
c2111 n1732__chipdriverout vss 119.514e-18
c2112 n1733__chipdriverout vss 126.924e-18
c2113 n731__i1__i14__net1 vss 37.9595e-18
c2114 n22__i5__i7__net44 vss 361.885e-18
c2115 n977__vddio vss 120.387e-18
c2116 n978__vddio vss 118.306e-18
c2117 n979__vddio vss 119.35e-18
c2118 n980__vddio vss 120.868e-18
c2119 n981__vddio vss 119.553e-18
c2120 n982__vddio vss 113.472e-18
c2121 n983__vddio vss 115.595e-18
c2122 n1126__vddio vss 76.9116e-18
c2123 n6__i5__r2 vss 19.9489e-18
c2124 n727__i1__i14__net1 vss 38.5537e-18
c2125 n1682__chipdriverout vss 133.582e-18
c2126 n1683__chipdriverout vss 108.863e-18
c2127 n1684__chipdriverout vss 120.567e-18
c2128 n1685__chipdriverout vss 108.308e-18
c2129 n1686__chipdriverout vss 74.9897e-18
c2130 n1687__chipdriverout vss 114.09e-18
c2131 n1688__chipdriverout vss 103.029e-18
c2132 n1689__chipdriverout vss 117.903e-18
c2133 n1690__chipdriverout vss 103.029e-18
c2134 n1691__chipdriverout vss 120.317e-18
c2135 n1692__chipdriverout vss 109.065e-18
c2136 n1693__chipdriverout vss 135.623e-18
c2137 n1694__chipdriverout vss 110.725e-18
c2138 n723__i1__i14__net1 vss 38.6692e-18
c2139 n956__vddio vss 102.77e-18
c2140 n957__vddio vss 134.625e-18
c2141 n958__vddio vss 103.421e-18
c2142 n959__vddio vss 104.699e-18
c2143 n960__vddio vss 103.421e-18
c2144 n961__vddio vss 129.794e-18
c2145 n962__vddio vss 99.6841e-18
c2146 n1127__vddio vss 77.551e-18
c2147 n719__i1__i14__net1 vss 40.7962e-18
c2148 n1643__chipdriverout vss 133.028e-18
c2149 n1644__chipdriverout vss 108.957e-18
c2150 n1645__chipdriverout vss 120.165e-18
c2151 n1646__chipdriverout vss 107.979e-18
c2152 n1647__chipdriverout vss 72.886e-18
c2153 n1648__chipdriverout vss 112.483e-18
c2154 n1649__chipdriverout vss 101.506e-18
c2155 n1650__chipdriverout vss 116.629e-18
c2156 n1651__chipdriverout vss 101.506e-18
c2157 n1652__chipdriverout vss 119.516e-18
c2158 n1653__chipdriverout vss 110.623e-18
c2159 n1654__chipdriverout vss 135.779e-18
c2160 n1655__chipdriverout vss 110.439e-18
c2161 n711__i1__i14__net1 vss 79.2638e-18
c2162 n13__shift vss 84.3559e-18
c2163 n935__vddio vss 138.965e-18
c2164 n936__vddio vss 137.305e-18
c2165 n937__vddio vss 138.023e-18
c2166 n938__vddio vss 139.524e-18
c2167 n939__vddio vss 119.029e-18
c2168 n940__vddio vss 113.372e-18
c2169 n941__vddio vss 115.074e-18
c2170 n1128__vddio vss 77.4736e-18
c2171 n22__i5__i7__i7__net1 vss 287.884e-18
c2172 n698__i1__i14__net1 vss 38.8985e-18
c2173 n15__i5__i6__net31 vss 24.4184e-18
c2174 n1604__chipdriverout vss 119.65e-18
c2175 n1605__chipdriverout vss 107.153e-18
c2176 n1606__chipdriverout vss 119.905e-18
c2177 n1607__chipdriverout vss 105.759e-18
c2178 n1608__chipdriverout vss 68.314e-18
c2179 n1609__chipdriverout vss 111.414e-18
c2180 n1610__chipdriverout vss 99.7454e-18
c2181 n1611__chipdriverout vss 114.93e-18
c2182 n1612__chipdriverout vss 99.7454e-18
c2183 n1613__chipdriverout vss 118.68e-18
c2184 n1614__chipdriverout vss 114.764e-18
c2185 n1615__chipdriverout vss 137.724e-18
c2186 n1616__chipdriverout vss 110.572e-18
c2187 n695__i1__i14__net1 vss 41.0098e-18
c2188 n914__vddio vss 104.945e-18
c2189 n915__vddio vss 136.649e-18
c2190 n916__vddio vss 105.552e-18
c2191 n917__vddio vss 106.831e-18
c2192 n918__vddio vss 104.148e-18
c2193 n919__vddio vss 129.79e-18
c2194 n920__vddio vss 98.8923e-18
c2195 n1129__vddio vss 54.64e-18
c2196 n6__i5__r1 vss 74.1545e-18
c2197 n681__i1__i14__net1 vss 39.6827e-18
c2198 n1564__chipdriverout vss 120.27e-18
c2199 n1565__chipdriverout vss 108.272e-18
c2200 n1566__chipdriverout vss 121.112e-18
c2201 n1567__chipdriverout vss 106.876e-18
c2202 n1568__chipdriverout vss 69.1306e-18
c2203 n1569__chipdriverout vss 112.191e-18
c2204 n1570__chipdriverout vss 100.929e-18
c2205 n1571__chipdriverout vss 116.247e-18
c2206 n1572__chipdriverout vss 100.929e-18
c2207 n1573__chipdriverout vss 121.922e-18
c2208 n1574__chipdriverout vss 108.724e-18
c2209 n1575__chipdriverout vss 139.392e-18
c2210 n1576__chipdriverout vss 107.833e-18
c2211 n16__i5__clk_buf vss 233.146e-18
c2212 n677__i1__i14__net1 vss 39.4476e-18
c2213 n869__vddio vss 122.675e-18
c2214 n872__vddio vss 120.795e-18
c2215 n873__vddio vss 121.652e-18
c2216 n876__vddio vss 123.171e-18
c2217 n877__vddio vss 120.448e-18
c2218 n880__vddio vss 113.689e-18
c2219 n881__vddio vss 113.414e-18
c2220 n1130__vddio vss 76.0467e-18
c2221 n665__i1__i14__net1 vss 39.5541e-18
c2222 n14__i5__i7__i6__net1 vss 141.038e-18
c2223 n1524__chipdriverout vss 104.103e-18
c2224 n1525__chipdriverout vss 108.278e-18
c2225 n1526__chipdriverout vss 137.525e-18
c2226 n1527__chipdriverout vss 106.874e-18
c2227 n1528__chipdriverout vss 69.1283e-18
c2228 n1529__chipdriverout vss 111.514e-18
c2229 n1530__chipdriverout vss 100.777e-18
c2230 n1531__chipdriverout vss 116.19e-18
c2231 n1532__chipdriverout vss 100.777e-18
c2232 n1533__chipdriverout vss 120.347e-18
c2233 n1534__chipdriverout vss 112.438e-18
c2234 n1535__chipdriverout vss 135.784e-18
c2235 n1536__chipdriverout vss 108.498e-18
c2236 n663__i1__i14__net1 vss 40.5792e-18
c2237 n12__i5__i7__net46 vss 72.277e-18
c2238 n9__i5__r0 vss 94.3446e-18
c2239 n49__vdd vss 281.149e-18
c2240 n862__vddio vss 122.785e-18
c2241 n863__vddio vss 120.486e-18
c2242 n864__vddio vss 121.375e-18
c2243 n865__vddio vss 122.888e-18
c2244 n866__vddio vss 120.224e-18
c2245 n867__vddio vss 114.359e-18
c2246 n868__vddio vss 116.243e-18
c2247 n1131__vddio vss 54.5586e-18
c2248 n655__i1__i14__net1 vss 48.1869e-18
c2249 n1445__chipdriverout vss 16.539e-18
c2250 n1449__chipdriverout vss 15.8803e-18
c2251 n1453__chipdriverout vss 17.764e-18
c2252 n1457__chipdriverout vss 15.3755e-18
c2253 n1461__chipdriverout vss 15.5803e-18
c2254 n1465__chipdriverout vss 15.3755e-18
c2255 n1469__chipdriverout vss 16.3643e-18
c2256 n642__i1__i14__net1 vss 76.1069e-18
c2257 n827__vddio vss 155.468e-18
c2258 n830__vddio vss 152.377e-18
c2259 n831__vddio vss 154.819e-18
c2260 n834__vddio vss 156.141e-18
c2261 n835__vddio vss 165.671e-18
c2262 n838__vddio vss 149.218e-18
c2263 n839__vddio vss 154.305e-18
c2264 n1132__vddio vss 85.0956e-18
c2265 n19__i5__i7__net51 vss 108.527e-18
c2266 n635__i1__i14__net1 vss 79.7196e-18
c2267 n18__i5__i7__net44 vss 248.421e-18
c2268 n1431__chipdriverout vss 14.9774e-18
c2269 n1432__chipdriverout vss 15.4231e-18
c2270 n1433__chipdriverout vss 15.1715e-18
c2271 n1434__chipdriverout vss 17.3292e-18
c2272 n1436__chipdriverout vss 15.1254e-18
c2273 n1437__chipdriverout vss 15.5662e-18
c2274 n1438__chipdriverout vss 15.3207e-18
c2275 n1440__chipdriverout vss 15.1254e-18
c2276 n1442__chipdriverout vss 15.641e-18
c2277 n5__i5__i7__net46 vss 100.092e-18
c2278 n1563__vddio vss 7.64793e-18
c2279 n627__i1__i14__net1 vss 48.4697e-18
c2280 n814__vddio vss 105.439e-18
c2281 n815__vddio vss 136.649e-18
c2282 n816__vddio vss 105.552e-18
c2283 n817__vddio vss 106.831e-18
c2284 n818__vddio vss 104.148e-18
c2285 n819__vddio vss 130.522e-18
c2286 n820__vddio vss 100.415e-18
c2287 n1133__vddio vss 54.1641e-18
c2288 n8__i5__i7__i6__net1 vss 168.367e-18
c2289 n623__i1__i14__net1 vss 40.7838e-18
c2290 n1391__chipdriverout vss 115.799e-18
c2291 n1392__chipdriverout vss 124.945e-18
c2292 n1393__chipdriverout vss 121.112e-18
c2293 n1394__chipdriverout vss 123.058e-18
c2294 n1395__chipdriverout vss 69.9668e-18
c2295 n1396__chipdriverout vss 112.342e-18
c2296 n1397__chipdriverout vss 100.929e-18
c2297 n1398__chipdriverout vss 132.471e-18
c2298 n1399__chipdriverout vss 100.929e-18
c2299 n1400__chipdriverout vss 119.824e-18
c2300 n1401__chipdriverout vss 115.558e-18
c2301 n1402__chipdriverout vss 138.329e-18
c2302 n1403__chipdriverout vss 111.267e-18
c2303 n615__i1__i14__net1 vss 47.4017e-18
c2304 n789__vddio vss 107.075e-18
c2305 n790__vddio vss 139.115e-18
c2306 n791__vddio vss 107.76e-18
c2307 n792__vddio vss 109.056e-18
c2308 n793__vddio vss 106.348e-18
c2309 n794__vddio vss 132.712e-18
c2310 n795__vddio vss 101.698e-18
c2311 n1134__vddio vss 56.2865e-18
c2312 n603__i1__i14__net1 vss 38.5305e-18
c2313 n1352__chipdriverout vss 121.493e-18
c2314 n1353__chipdriverout vss 125.411e-18
c2315 n1354__chipdriverout vss 122.13e-18
c2316 n1355__chipdriverout vss 124.203e-18
c2317 n1356__chipdriverout vss 88.2084e-18
c2318 n1357__chipdriverout vss 90.9757e-18
c2319 n1358__chipdriverout vss 118.715e-18
c2320 n1359__chipdriverout vss 134.738e-18
c2321 n1360__chipdriverout vss 118.939e-18
c2322 n1361__chipdriverout vss 107.267e-18
c2323 n1362__chipdriverout vss 129.127e-18
c2324 n1363__chipdriverout vss 125.334e-18
c2325 n1364__chipdriverout vss 126.885e-18
c2326 n11__i5__i7__net47 vss 296.682e-18
c2327 n17__i5__i7__net51 vss 33.8443e-18
c2328 n599__i1__i14__net1 vss 40.3163e-18
c2329 n51__vdd vss 194.527e-18
c2330 n768__vddio vss 105.376e-18
c2331 n769__vddio vss 137.238e-18
c2332 n770__vddio vss 105.988e-18
c2333 n771__vddio vss 107.272e-18
c2334 n772__vddio vss 104.636e-18
c2335 n773__vddio vss 129.156e-18
c2336 n774__vddio vss 97.5405e-18
c2337 n1135__vddio vss 76.5875e-18
c2338 n586__i1__i14__net1 vss 38.2845e-18
c2339 n1313__chipdriverout vss 120.937e-18
c2340 n1314__chipdriverout vss 108.756e-18
c2341 n1315__chipdriverout vss 121.766e-18
c2342 n1316__chipdriverout vss 107.354e-18
c2343 n1317__chipdriverout vss 69.3251e-18
c2344 n1318__chipdriverout vss 112.343e-18
c2345 n1319__chipdriverout vss 101.436e-18
c2346 n1320__chipdriverout vss 116.984e-18
c2347 n1321__chipdriverout vss 101.436e-18
c2348 n1322__chipdriverout vss 121.787e-18
c2349 n1323__chipdriverout vss 112.705e-18
c2350 n1324__chipdriverout vss 142.619e-18
c2351 n1325__chipdriverout vss 109.833e-18
c2352 n8__i5__i7__net44 vss 339.356e-18
c2353 n583__i1__i14__net1 vss 39.1282e-18
c2354 n747__vddio vss 121.168e-18
c2355 n748__vddio vss 152.874e-18
c2356 n749__vddio vss 121.815e-18
c2357 n750__vddio vss 123.075e-18
c2358 n751__vddio vss 102.72e-18
c2359 n752__vddio vss 129.037e-18
c2360 n753__vddio vss 98.5162e-18
c2361 n1136__vddio vss 53.8535e-18
c2362 n14__i5__i7__i5__net1 vss 190.758e-18
c2363 n14__i5__i7__i4__net1 vss 122.585e-18
c2364 n575__i1__i14__net1 vss 79.8378e-18
c2365 n1274__chipdriverout vss 101.674e-18
c2366 n1275__chipdriverout vss 106.192e-18
c2367 n1276__chipdriverout vss 119.143e-18
c2368 n1277__chipdriverout vss 120.984e-18
c2369 n1278__chipdriverout vss 90.9884e-18
c2370 n1279__chipdriverout vss 89.8563e-18
c2371 n1280__chipdriverout vss 117.703e-18
c2372 n1281__chipdriverout vss 133.008e-18
c2373 n1282__chipdriverout vss 117.917e-18
c2374 n1283__chipdriverout vss 103.332e-18
c2375 n1284__chipdriverout vss 125.702e-18
c2376 n1285__chipdriverout vss 118.738e-18
c2377 n1286__chipdriverout vss 126.27e-18
c2378 n13__i5__i7__net51 vss 174.377e-18
c2379 n1567__vddio vss 6.80518e-18
c2380 n567__i1__i14__net1 vss 35.7718e-18
c2381 n726__vddio vss 120.494e-18
c2382 n727__vddio vss 118.39e-18
c2383 n728__vddio vss 119.371e-18
c2384 n729__vddio vss 120.886e-18
c2385 n730__vddio vss 119.574e-18
c2386 n731__vddio vss 113.506e-18
c2387 n732__vddio vss 115.953e-18
c2388 n1137__vddio vss 84.1058e-18
c2389 n559__i1__i14__net1 vss 38.5342e-18
c2390 n1235__chipdriverout vss 144.72e-18
c2391 n1236__chipdriverout vss 108.334e-18
c2392 n1237__chipdriverout vss 120.024e-18
c2393 n1238__chipdriverout vss 107.727e-18
c2394 n1239__chipdriverout vss 75.3564e-18
c2395 n1240__chipdriverout vss 114.474e-18
c2396 n1241__chipdriverout vss 103.295e-18
c2397 n1242__chipdriverout vss 118.126e-18
c2398 n1243__chipdriverout vss 103.295e-18
c2399 n1244__chipdriverout vss 120.821e-18
c2400 n1245__chipdriverout vss 109.528e-18
c2401 n1246__chipdriverout vss 136.058e-18
c2402 n1247__chipdriverout vss 111.343e-18
c2403 n551__i1__i14__net1 vss 30.8485e-18
c2404 n19__i5__i7__xor2 vss 149.548e-18
c2405 n18__i5__i7__xor1 vss 103.065e-18
c2406 n705__vddio vss 123.251e-18
c2407 n706__vddio vss 121.299e-18
c2408 n707__vddio vss 122.08e-18
c2409 n708__vddio vss 123.624e-18
c2410 n709__vddio vss 122.283e-18
c2411 n710__vddio vss 116.289e-18
c2412 n711__vddio vss 118.221e-18
c2413 n1138__vddio vss 55.2752e-18
c2414 n539__i1__i14__net1 vss 39.2702e-18
c2415 n6__i5__i7__net47 vss 187.501e-18
c2416 n5__i5__i7__net44 vss 268.163e-18
c2417 n1196__chipdriverout vss 140.665e-18
c2418 n1197__chipdriverout vss 126.651e-18
c2419 n1198__chipdriverout vss 122.312e-18
c2420 n1199__chipdriverout vss 125.795e-18
c2421 n1200__chipdriverout vss 95.9063e-18
c2422 n1201__chipdriverout vss 93.371e-18
c2423 n1202__chipdriverout vss 122.147e-18
c2424 n1203__chipdriverout vss 137.709e-18
c2425 n1204__chipdriverout vss 122.371e-18
c2426 n1205__chipdriverout vss 107.435e-18
c2427 n1206__chipdriverout vss 128.326e-18
c2428 n1207__chipdriverout vss 122.775e-18
c2429 n1208__chipdriverout vss 129.877e-18
c2430 n535__i1__i14__net1 vss 36.278e-18
c2431 n11__i5__i7__i5__net1 vss 196.638e-18
c2432 n11__i5__i7__i4__net1 vss 262.056e-18
c2433 n53__vdd vss 148.973e-18
c2434 n670__vddio vss 122.465e-18
c2435 n673__vddio vss 120.692e-18
c2436 n674__vddio vss 121.396e-18
c2437 n677__vddio vss 122.94e-18
c2438 n678__vddio vss 121.598e-18
c2439 n681__vddio vss 115.729e-18
c2440 n682__vddio vss 117.565e-18
c2441 n1139__vddio vss 55.3589e-18
c2442 n521__i1__i14__net1 vss 37.258e-18
c2443 n1157__chipdriverout vss 105.101e-18
c2444 n1158__chipdriverout vss 125.432e-18
c2445 n1159__chipdriverout vss 138.925e-18
c2446 n1160__chipdriverout vss 124.215e-18
c2447 n1161__chipdriverout vss 94.838e-18
c2448 n1162__chipdriverout vss 92.5849e-18
c2449 n1163__chipdriverout vss 121.603e-18
c2450 n1164__chipdriverout vss 137.301e-18
c2451 n1165__chipdriverout vss 121.817e-18
c2452 n1166__chipdriverout vss 106.929e-18
c2453 n1167__chipdriverout vss 128.724e-18
c2454 n1168__chipdriverout vss 122.413e-18
c2455 n1169__chipdriverout vss 129.388e-18
c2456 n519__i1__i14__net1 vss 36.1122e-18
c2457 n663__vddio vss 118.914e-18
c2458 n664__vddio vss 116.923e-18
c2459 n665__vddio vss 117.898e-18
c2460 n666__vddio vss 119.403e-18
c2461 n667__vddio vss 118.1e-18
c2462 n668__vddio vss 111.682e-18
c2463 n669__vddio vss 112.801e-18
c2464 n1140__vddio vss 53.651e-18
c2465 n511__i1__i14__net1 vss 37.2878e-18
c2466 n17__i5__i7__xor2 vss 21.528e-18
c2467 n17__i5__i7__xor1 vss 74.4991e-18
c2468 n1092__chipdriverout vss 101.44e-18
c2469 n1095__chipdriverout vss 121.842e-18
c2470 n1096__chipdriverout vss 135.15e-18
c2471 n1099__chipdriverout vss 120.673e-18
c2472 n1100__chipdriverout vss 90.9463e-18
c2473 n1103__chipdriverout vss 89.4947e-18
c2474 n1104__chipdriverout vss 118.155e-18
c2475 n1107__chipdriverout vss 133.484e-18
c2476 n1108__chipdriverout vss 118.363e-18
c2477 n1111__chipdriverout vss 106.547e-18
c2478 n1112__chipdriverout vss 128.812e-18
c2479 n1115__chipdriverout vss 123.585e-18
c2480 n1116__chipdriverout vss 122.508e-18
c2481 n1571__vddio vss 6.98695e-18
c2482 n503__i1__i14__net1 vss 36.1015e-18
c2483 n632__vddio vss 119.695e-18
c2484 n633__vddio vss 117.55e-18
c2485 n634__vddio vss 118.571e-18
c2486 n635__vddio vss 120.076e-18
c2487 n636__vddio vss 118.774e-18
c2488 n637__vddio vss 111.417e-18
c2489 n638__vddio vss 111.438e-18
c2490 n1141__vddio vss 81.1744e-18
c2491 n491__i1__i14__net1 vss 38.0258e-18
c2492 n1079__chipdriverout vss 102.122e-18
c2493 n1080__chipdriverout vss 121.79e-18
c2494 n1081__chipdriverout vss 134.952e-18
c2495 n1082__chipdriverout vss 120.621e-18
c2496 n1083__chipdriverout vss 90.7444e-18
c2497 n1084__chipdriverout vss 89.8977e-18
c2498 n1085__chipdriverout vss 118.376e-18
c2499 n1086__chipdriverout vss 133.55e-18
c2500 n1087__chipdriverout vss 118.594e-18
c2501 n1088__chipdriverout vss 105.302e-18
c2502 n1089__chipdriverout vss 129.109e-18
c2503 n1090__chipdriverout vss 123.412e-18
c2504 n1091__chipdriverout vss 128.9e-18
c2505 n487__i1__i14__net1 vss 35.3358e-18
c2506 n597__vddio vss 123.188e-18
c2507 n600__vddio vss 121.131e-18
c2508 n601__vddio vss 121.955e-18
c2509 n604__vddio vss 123.499e-18
c2510 n605__vddio vss 122.157e-18
c2511 n608__vddio vss 116.117e-18
c2512 n609__vddio vss 117.97e-18
c2513 n1142__vddio vss 77.9818e-18
c2514 n475__i1__i14__net1 vss 38.0774e-18
c2515 n1040__chipdriverout vss 133.881e-18
c2516 n1041__chipdriverout vss 125.929e-18
c2517 n1042__chipdriverout vss 122.321e-18
c2518 n1043__chipdriverout vss 124.102e-18
c2519 n1044__chipdriverout vss 93.872e-18
c2520 n1045__chipdriverout vss 92.992e-18
c2521 n1046__chipdriverout vss 121.933e-18
c2522 n1047__chipdriverout vss 137.447e-18
c2523 n1048__chipdriverout vss 122.151e-18
c2524 n1049__chipdriverout vss 107.205e-18
c2525 n1050__chipdriverout vss 128.159e-18
c2526 n1051__chipdriverout vss 122.476e-18
c2527 n1052__chipdriverout vss 130.158e-18
c2528 n469__i1__i14__net1 vss 35.9087e-18
c2529 n55__vdd vss 271.166e-18
c2530 n590__vddio vss 121.268e-18
c2531 n591__vddio vss 119.273e-18
c2532 n592__vddio vss 120.163e-18
c2533 n593__vddio vss 121.698e-18
c2534 n594__vddio vss 120.365e-18
c2535 n595__vddio vss 114.356e-18
c2536 n596__vddio vss 116.359e-18
c2537 n1143__vddio vss 77.6306e-18
c2538 n463__i1__i14__net1 vss 40.0483e-18
c2539 n975__chipdriverout vss 114.98e-18
c2540 n978__chipdriverout vss 124.562e-18
c2541 n979__chipdriverout vss 138.178e-18
c2542 n982__chipdriverout vss 125.276e-18
c2543 n983__chipdriverout vss 95.4768e-18
c2544 n986__chipdriverout vss 91.509e-18
c2545 n987__chipdriverout vss 120.713e-18
c2546 n990__chipdriverout vss 136.386e-18
c2547 n991__chipdriverout vss 120.918e-18
c2548 n994__chipdriverout vss 106.155e-18
c2549 n995__chipdriverout vss 127.667e-18
c2550 n998__chipdriverout vss 121.585e-18
c2551 n999__chipdriverout vss 133.768e-18
c2552 n455__i1__i14__net1 vss 38.6324e-18
c2553 n13__i5__i7__y3out vss 293.652e-18
c2554 n545__vddio vss 121.132e-18
c2555 n548__vddio vss 119.391e-18
c2556 n549__vddio vss 120.129e-18
c2557 n552__vddio vss 121.653e-18
c2558 n553__vddio vss 120.332e-18
c2559 n556__vddio vss 114.516e-18
c2560 n557__vddio vss 116.654e-18
c2561 n1144__vddio vss 54.5193e-18
c2562 n11__i5__i7__x3out vss 80.9887e-18
c2563 n12__i5__i7__x0out vss 60.5701e-18
c2564 n445__i1__i14__net1 vss 38.7763e-18
c2565 n962__chipdriverout vss 122.498e-18
c2566 n963__chipdriverout vss 125.394e-18
c2567 n964__chipdriverout vss 136.996e-18
c2568 n965__chipdriverout vss 124.271e-18
c2569 n966__chipdriverout vss 94.7162e-18
c2570 n967__chipdriverout vss 91.4802e-18
c2571 n968__chipdriverout vss 120.17e-18
c2572 n969__chipdriverout vss 135.551e-18
c2573 n970__chipdriverout vss 120.378e-18
c2574 n971__chipdriverout vss 105.54e-18
c2575 n972__chipdriverout vss 127.539e-18
c2576 n973__chipdriverout vss 122.617e-18
c2577 n974__chipdriverout vss 128.271e-18
c2578 n1575__vddio vss 6.1597e-18
c2579 n439__i1__i14__net1 vss 35.4787e-18
c2580 n538__vddio vss 123.001e-18
c2581 n539__vddio vss 121.303e-18
c2582 n540__vddio vss 121.965e-18
c2583 n541__vddio vss 123.515e-18
c2584 n542__vddio vss 122.168e-18
c2585 n543__vddio vss 115.725e-18
c2586 n544__vddio vss 116.299e-18
c2587 n1145__vddio vss 77.9858e-18
c2588 n429__i1__i14__net1 vss 37.7459e-18
c2589 n923__chipdriverout vss 103.963e-18
c2590 n924__chipdriverout vss 124.355e-18
c2591 n925__chipdriverout vss 137.389e-18
c2592 n926__chipdriverout vss 123.076e-18
c2593 n927__chipdriverout vss 92.993e-18
c2594 n928__chipdriverout vss 93.6502e-18
c2595 n929__chipdriverout vss 122.146e-18
c2596 n930__chipdriverout vss 137.712e-18
c2597 n931__chipdriverout vss 122.353e-18
c2598 n932__chipdriverout vss 111.076e-18
c2599 n933__chipdriverout vss 131.933e-18
c2600 n934__chipdriverout vss 125.626e-18
c2601 n935__chipdriverout vss 125.181e-18
c2602 n419__i1__i14__net1 vss 36.5455e-18
c2603 n10__i5__i7__xor2 vss 211.968e-18
c2604 n10__i5__i7__xor1 vss 193.193e-18
c2605 n517__vddio vss 119.401e-18
c2606 n518__vddio vss 133.747e-18
c2607 n519__vddio vss 118.427e-18
c2608 n520__vddio vss 119.944e-18
c2609 n521__vddio vss 118.628e-18
c2610 n522__vddio vss 111.832e-18
c2611 n523__vddio vss 111.872e-18
c2612 n1146__vddio vss 53.6527e-18
c2613 n411__i1__i14__net1 vss 38.1463e-18
c2614 n892__chipdriverout vss 102.276e-18
c2615 n893__chipdriverout vss 106.737e-18
c2616 n894__chipdriverout vss 119.191e-18
c2617 n895__chipdriverout vss 105.44e-18
c2618 n896__chipdriverout vss 73.1321e-18
c2619 n873__chipdriverout vss 90.993e-18
c2620 n874__chipdriverout vss 103.112e-18
c2621 n875__chipdriverout vss 118.173e-18
c2622 n876__chipdriverout vss 103.112e-18
c2623 n877__chipdriverout vss 121.417e-18
c2624 n878__chipdriverout vss 113.576e-18
c2625 n879__chipdriverout vss 123.758e-18
c2626 n880__chipdriverout vss 109.227e-18
c2627 n403__i1__i14__net1 vss 37.2934e-18
c2628 n57__vdd vss 225.113e-18
c2629 n496__vddio vss 101.657e-18
c2630 n497__vddio vss 133.529e-18
c2631 n498__vddio vss 102.367e-18
c2632 n499__vddio vss 103.63e-18
c2633 n500__vddio vss 102.367e-18
c2634 n501__vddio vss 128.739e-18
c2635 n502__vddio vss 98.9583e-18
c2636 n1147__vddio vss 81.3102e-18
c2637 n398__i1__i14__net1 vss 36.4032e-18
c2638 n845__chipdriverout vss 123.249e-18
c2639 n846__chipdriverout vss 125.71e-18
c2640 n847__chipdriverout vss 137.534e-18
c2641 n848__chipdriverout vss 124.537e-18
c2642 n849__chipdriverout vss 95.5258e-18
c2643 n850__chipdriverout vss 90.5008e-18
c2644 n851__chipdriverout vss 118.324e-18
c2645 n852__chipdriverout vss 133.522e-18
c2646 n853__chipdriverout vss 118.532e-18
c2647 n854__chipdriverout vss 103.723e-18
c2648 n855__chipdriverout vss 124.268e-18
c2649 n856__chipdriverout vss 118.67e-18
c2650 n857__chipdriverout vss 131.246e-18
c2651 n11__i5__i7__x2out vss 88.0815e-18
c2652 n387__i1__i14__net1 vss 37.5233e-18
c2653 n12__i5__i7__x1out vss 87.2745e-18
c2654 n475__vddio vss 103.821e-18
c2655 n476__vddio vss 135.649e-18
c2656 n477__vddio vss 104.445e-18
c2657 n478__vddio vss 105.732e-18
c2658 n479__vddio vss 104.445e-18
c2659 n480__vddio vss 130.776e-18
c2660 n481__vddio vss 100.988e-18
c2661 n1148__vddio vss 81.6743e-18
c2662 n383__i1__i14__net1 vss 41.8664e-18
c2663 n11__i5__i7__y3out vss 198.323e-18
c2664 n806__chipdriverout vss 107.088e-18
c2665 n807__chipdriverout vss 121.614e-18
c2666 n808__chipdriverout vss 136.469e-18
c2667 n809__chipdriverout vss 121.816e-18
c2668 n810__chipdriverout vss 95.2481e-18
c2669 n811__chipdriverout vss 92.3842e-18
c2670 n812__chipdriverout vss 120.369e-18
c2671 n813__chipdriverout vss 135.77e-18
c2672 n814__chipdriverout vss 120.576e-18
c2673 n815__chipdriverout vss 105.724e-18
c2674 n816__chipdriverout vss 127.316e-18
c2675 n817__chipdriverout vss 120.877e-18
c2676 n818__chipdriverout vss 128.407e-18
c2677 n1579__vddio vss 7.07332e-18
c2678 n371__i1__i14__net1 vss 46.8168e-18
c2679 n34__reset vss 185.744e-18
c2680 n33__reset vss 139.783e-18
c2681 n434__vddio vss 122.945e-18
c2682 n437__vddio vss 121.175e-18
c2683 n438__vddio vss 121.878e-18
c2684 n441__vddio vss 123.424e-18
c2685 n442__vddio vss 122.08e-18
c2686 n445__vddio vss 116.213e-18
c2687 n446__vddio vss 118.048e-18
c2688 n1149__vddio vss 79.2554e-18
c2689 n367__i1__i14__net1 vss 29.2467e-18
c2690 n767__chipdriverout vss 141.515e-18
c2691 n768__chipdriverout vss 112.457e-18
c2692 n769__chipdriverout vss 123.407e-18
c2693 n770__chipdriverout vss 110.863e-18
c2694 n771__chipdriverout vss 75.9396e-18
c2695 n772__chipdriverout vss 117.093e-18
c2696 n773__chipdriverout vss 105.828e-18
c2697 n774__chipdriverout vss 120.842e-18
c2698 n775__chipdriverout vss 105.828e-18
c2699 n776__chipdriverout vss 123.384e-18
c2700 n777__chipdriverout vss 111.988e-18
c2701 n778__chipdriverout vss 138.763e-18
c2702 n779__chipdriverout vss 113.26e-18
c2703 n355__i1__i14__net1 vss 37.1091e-18
c2704 n410__vddio vss 104.409e-18
c2705 n411__vddio vss 136.27e-18
c2706 n414__vddio vss 104.924e-18
c2707 n415__vddio vss 106.225e-18
c2708 n418__vddio vss 104.924e-18
c2709 n419__vddio vss 131.253e-18
c2710 n422__vddio vss 100.317e-18
c2711 n1150__vddio vss 54.6244e-18
c2712 n351__i1__i14__net1 vss 35.9405e-18
c2713 n728__chipdriverout vss 104.403e-18
c2714 n729__chipdriverout vss 124.551e-18
c2715 n730__chipdriverout vss 138.057e-18
c2716 n731__chipdriverout vss 123.343e-18
c2717 n732__chipdriverout vss 92.8697e-18
c2718 n733__chipdriverout vss 92.7335e-18
c2719 n734__chipdriverout vss 120.867e-18
c2720 n735__chipdriverout vss 136.391e-18
c2721 n736__chipdriverout vss 121.075e-18
c2722 n737__chipdriverout vss 108.471e-18
c2723 n738__chipdriverout vss 141.747e-18
c2724 n739__chipdriverout vss 125.993e-18
c2725 n740__chipdriverout vss 125.686e-18
c2726 n339__i1__i14__net1 vss 36.4865e-18
c2727 n389__vddio vss 102.658e-18
c2728 n390__vddio vss 134.605e-18
c2729 n393__vddio vss 103.353e-18
c2730 n394__vddio vss 104.628e-18
c2731 n397__vddio vss 103.353e-18
c2732 n398__vddio vss 127.792e-18
c2733 n401__vddio vss 96.2617e-18
c2734 n1151__vddio vss 75.7307e-18
c2735 n68__i5__clk4 vss 305.937e-18
c2736 n30__i5__i7__i1__net1 vss 299.91e-18
c2737 n64__i5__clk4 vss 280.164e-18
c2738 n30__i5__i7__i0__net1 vss 306.868e-18
c2739 n331__i1__i14__net1 vss 37.4787e-18
c2740 n689__chipdriverout vss 102.285e-18
c2741 n690__chipdriverout vss 122.687e-18
c2742 n691__chipdriverout vss 136.009e-18
c2743 n692__chipdriverout vss 121.51e-18
c2744 n693__chipdriverout vss 91.7932e-18
c2745 n694__chipdriverout vss 91.3061e-18
c2746 n695__chipdriverout vss 119.104e-18
c2747 n696__chipdriverout vss 134.408e-18
c2748 n697__chipdriverout vss 119.311e-18
c2749 n698__chipdriverout vss 107.041e-18
c2750 n699__chipdriverout vss 139.461e-18
c2751 n700__chipdriverout vss 124.869e-18
c2752 n701__chipdriverout vss 124.203e-18
c2753 n323__i1__i14__net1 vss 34.7167e-18
c2754 n367__vddio vss 121.597e-18
c2755 n370__vddio vss 119.431e-18
c2756 n371__vddio vss 120.406e-18
c2757 n374__vddio vss 121.934e-18
c2758 n375__vddio vss 120.609e-18
c2759 n378__vddio vss 114.364e-18
c2760 n379__vddio vss 116.348e-18
c2761 n1152__vddio vss 53.8983e-18
c2762 n5__y3 vss 29.7406e-18
c2763 n318__i1__i14__net1 vss 35.4603e-18
c2764 n650__chipdriverout vss 116.296e-18
c2765 n651__chipdriverout vss 125.378e-18
c2766 n652__chipdriverout vss 121.194e-18
c2767 n653__chipdriverout vss 107.158e-18
c2768 n654__chipdriverout vss 94.052e-18
c2769 n655__chipdriverout vss 91.9456e-18
c2770 n656__chipdriverout vss 104.506e-18
c2771 n657__chipdriverout vss 119.557e-18
c2772 n658__chipdriverout vss 120.466e-18
c2773 n659__chipdriverout vss 105.79e-18
c2774 n660__chipdriverout vss 127.015e-18
c2775 n661__chipdriverout vss 121.057e-18
c2776 n662__chipdriverout vss 133.806e-18
c2777 n311__i1__i14__net1 vss 34.928e-18
c2778 n9__i5__i7__x2out vss 61.8294e-18
c2779 n346__vddio vss 121.154e-18
c2780 n349__vddio vss 119.439e-18
c2781 n350__vddio vss 120.117e-18
c2782 n353__vddio vss 121.639e-18
c2783 n354__vddio vss 120.319e-18
c2784 n357__vddio vss 114.566e-18
c2785 n358__vddio vss 116.338e-18
c2786 n1153__vddio vss 77.0519e-18
c2787 n30__reset vss 357.085e-18
c2788 n28__reset vss 326.145e-18
c2789 n298__i1__i14__net1 vss 37.9068e-18
c2790 n611__chipdriverout vss 130.235e-18
c2791 n612__chipdriverout vss 108.471e-18
c2792 n613__chipdriverout vss 121.564e-18
c2793 n614__chipdriverout vss 109.007e-18
c2794 n615__chipdriverout vss 76.6437e-18
c2795 n616__chipdriverout vss 114.739e-18
c2796 n617__chipdriverout vss 104.078e-18
c2797 n618__chipdriverout vss 119.163e-18
c2798 n619__chipdriverout vss 104.078e-18
c2799 n620__chipdriverout vss 121.413e-18
c2800 n621__chipdriverout vss 110.364e-18
c2801 n622__chipdriverout vss 136.895e-18
c2802 n623__chipdriverout vss 111.53e-18
c2803 n291__i1__i14__net1 vss 37.8101e-18
c2804 n339__vddio vss 103.469e-18
c2805 n340__vddio vss 135.525e-18
c2806 n341__vddio vss 104.167e-18
c2807 n342__vddio vss 105.449e-18
c2808 n343__vddio vss 104.167e-18
c2809 n344__vddio vss 130.653e-18
c2810 n345__vddio vss 100.405e-18
c2811 n1154__vddio vss 54.3882e-18
c2812 n283__i1__i14__net1 vss 39.3495e-18
c2813 n547__chipdriverout vss 139.792e-18
c2814 n548__chipdriverout vss 109.939e-18
c2815 n551__chipdriverout vss 121.217e-18
c2816 n552__chipdriverout vss 108.633e-18
c2817 n555__chipdriverout vss 77.0488e-18
c2818 n556__chipdriverout vss 115.136e-18
c2819 n559__chipdriverout vss 103.979e-18
c2820 n560__chipdriverout vss 118.98e-18
c2821 n563__chipdriverout vss 103.979e-18
c2822 n564__chipdriverout vss 121.377e-18
c2823 n567__chipdriverout vss 110.013e-18
c2824 n568__chipdriverout vss 136.761e-18
c2825 n571__chipdriverout vss 111.499e-18
c2826 n277__i1__i14__net1 vss 38.0348e-18
c2827 n304__vddio vss 121.472e-18
c2828 n307__vddio vss 119.248e-18
c2829 n308__vddio vss 120.292e-18
c2830 n311__vddio vss 121.819e-18
c2831 n312__vddio vss 120.494e-18
c2832 n315__vddio vss 114.319e-18
c2833 n316__vddio vss 116.481e-18
c2834 n1155__vddio vss 77.963e-18
c2835 n267__i1__i14__net1 vss 28.5852e-18
c2836 n29__i5__i7__i1__net1 vss 242.756e-18
c2837 n29__i5__i7__i0__net1 vss 436.814e-18
c2838 n508__chipdriverout vss 120.301e-18
c2839 n509__chipdriverout vss 108.355e-18
c2840 n512__chipdriverout vss 121.194e-18
c2841 n513__chipdriverout vss 106.951e-18
c2842 n516__chipdriverout vss 75.7415e-18
c2843 n517__chipdriverout vss 115.079e-18
c2844 n520__chipdriverout vss 104.407e-18
c2845 n521__chipdriverout vss 119.374e-18
c2846 n524__chipdriverout vss 104.408e-18
c2847 n525__chipdriverout vss 121.748e-18
c2848 n528__chipdriverout vss 111.412e-18
c2849 n529__chipdriverout vss 137.115e-18
c2850 n532__chipdriverout vss 111.738e-18
c2851 n263__i1__i14__net1 vss 38.005e-18
c2852 n297__vddio vss 122.309e-18
c2853 n298__vddio vss 120.237e-18
c2854 n299__vddio vss 121.14e-18
c2855 n300__vddio vss 122.676e-18
c2856 n301__vddio vss 121.343e-18
c2857 n302__vddio vss 114.785e-18
c2858 n303__vddio vss 116.104e-18
c2859 n1156__vddio vss 55.142e-18
c2860 n250__i1__i14__net1 vss 35.9418e-18
c2861 n7__y2 vss 23.082e-18
c2862 n494__chipdriverout vss 124.09e-18
c2863 n495__chipdriverout vss 108.857e-18
c2864 n496__chipdriverout vss 121.646e-18
c2865 n497__chipdriverout vss 107.452e-18
c2866 n498__chipdriverout vss 74.4099e-18
c2867 n499__chipdriverout vss 115.659e-18
c2868 n500__chipdriverout vss 104.977e-18
c2869 n501__chipdriverout vss 120.014e-18
c2870 n502__chipdriverout vss 104.977e-18
c2871 n503__chipdriverout vss 125.356e-18
c2872 n504__chipdriverout vss 116.083e-18
c2873 n505__chipdriverout vss 142.653e-18
c2874 n506__chipdriverout vss 109.951e-18
c2875 n1587__vddio vss 7.2337e-18
c2876 n247__i1__i14__net1 vss 37.9538e-18
c2877 n6__i5__i7__y1out vss 108.913e-18
c2878 n6__i5__i7__x1out vss 38.7731e-18
c2879 n266__vddio vss 102.813e-18
c2880 n267__vddio vss 134.668e-18
c2881 n268__vddio vss 103.423e-18
c2882 n269__vddio vss 104.7e-18
c2883 n270__vddio vss 103.423e-18
c2884 n271__vddio vss 128.078e-18
c2885 n272__vddio vss 96.5806e-18
c2886 n1157__vddio vss 54.1009e-18
c2887 n235__i1__i14__net1 vss 43.5544e-18
c2888 n23__reset vss 358.1e-18
c2889 n22__reset vss 362.016e-18
c2890 n455__chipdriverout vss 119.47e-18
c2891 n456__chipdriverout vss 107.194e-18
c2892 n457__chipdriverout vss 120.076e-18
c2893 n458__chipdriverout vss 105.802e-18
c2894 n459__chipdriverout vss 73.3916e-18
c2895 n460__chipdriverout vss 114.127e-18
c2896 n461__chipdriverout vss 103.38e-18
c2897 n462__chipdriverout vss 118.309e-18
c2898 n463__chipdriverout vss 103.38e-18
c2899 n464__chipdriverout vss 122.432e-18
c2900 n465__chipdriverout vss 114.109e-18
c2901 n466__chipdriverout vss 140.707e-18
c2902 n467__chipdriverout vss 108.349e-18
c2903 n231__i1__i14__net1 vss 38.7884e-18
c2904 n231__vddio vss 119.378e-18
c2905 n234__vddio vss 117.578e-18
c2906 n235__vddio vss 118.409e-18
c2907 n238__vddio vss 119.914e-18
c2908 n239__vddio vss 118.612e-18
c2909 n242__vddio vss 112.79e-18
c2910 n243__vddio vss 114.592e-18
c2911 n1158__vddio vss 76.525e-18
c2912 n223__i1__i14__net1 vss 37.6298e-18
c2913 n416__chipdriverout vss 130.631e-18
c2914 n417__chipdriverout vss 107.99e-18
c2915 n418__chipdriverout vss 118.889e-18
c2916 n419__chipdriverout vss 104.828e-18
c2917 n420__chipdriverout vss 74.146e-18
c2918 n421__chipdriverout vss 113.263e-18
c2919 n422__chipdriverout vss 102.348e-18
c2920 n423__chipdriverout vss 117.107e-18
c2921 n424__chipdriverout vss 102.348e-18
c2922 n425__chipdriverout vss 119.584e-18
c2923 n426__chipdriverout vss 109.235e-18
c2924 n427__chipdriverout vss 134.728e-18
c2925 n428__chipdriverout vss 109.926e-18
c2926 n215__i1__i14__net1 vss 37.7248e-18
c2927 n63__vdd vss 200.09e-18
c2928 n224__vddio vss 103.96e-18
c2929 n225__vddio vss 135.774e-18
c2930 n226__vddio vss 104.596e-18
c2931 n227__vddio vss 105.883e-18
c2932 n228__vddio vss 104.596e-18
c2933 n229__vddio vss 130.902e-18
c2934 n230__vddio vss 100.834e-18
c2935 n1159__vddio vss 77.5206e-18
c2936 n206__i1__i14__net1 vss 38.7704e-18
c2937 n377__chipdriverout vss 114.444e-18
c2938 n378__chipdriverout vss 108.345e-18
c2939 n379__chipdriverout vss 121.285e-18
c2940 n380__chipdriverout vss 108.845e-18
c2941 n381__chipdriverout vss 76.7588e-18
c2942 n382__chipdriverout vss 114.844e-18
c2943 n383__chipdriverout vss 104.429e-18
c2944 n384__chipdriverout vss 119.499e-18
c2945 n385__chipdriverout vss 104.429e-18
c2946 n386__chipdriverout vss 121.777e-18
c2947 n387__chipdriverout vss 111.371e-18
c2948 n388__chipdriverout vss 137.259e-18
c2949 n389__chipdriverout vss 111.768e-18
c2950 n24__i5__i7__i1__net1 vss 397.427e-18
c2951 n24__i5__i7__i0__net1 vss 423.127e-18
c2952 n193__i1__i14__net1 vss 39.8197e-18
c2953 n193__vddio vss 103.436e-18
c2954 n194__vddio vss 135.445e-18
c2955 n195__vddio vss 104.155e-18
c2956 n196__vddio vss 105.436e-18
c2957 n197__vddio vss 104.155e-18
c2958 n198__vddio vss 130.518e-18
c2959 n199__vddio vss 100.665e-18
c2960 n1160__vddio vss 83.5362e-18
c2961 n191__i1__i14__net1 vss 36.2984e-18
c2962 n338__chipdriverout vss 142.625e-18
c2963 n339__chipdriverout vss 110.552e-18
c2964 n340__chipdriverout vss 121.326e-18
c2965 n341__chipdriverout vss 108.573e-18
c2966 n342__chipdriverout vss 92.4213e-18
c2967 n343__chipdriverout vss 114.236e-18
c2968 n344__chipdriverout vss 104.287e-18
c2969 n345__chipdriverout vss 119.329e-18
c2970 n346__chipdriverout vss 104.287e-18
c2971 n347__chipdriverout vss 139.36e-18
c2972 n348__chipdriverout vss 124.869e-18
c2973 n349__chipdriverout vss 138.008e-18
c2974 n350__chipdriverout vss 112.29e-18
c2975 n5__y1 vss 24.0249e-18
c2976 n5__x1 vss 23.8347e-18
c2977 n183__i1__i14__net1 vss 81.5508e-18
c2978 n172__vddio vss 103.319e-18
c2979 n173__vddio vss 135.32e-18
c2980 n174__vddio vss 119.873e-18
c2981 n175__vddio vss 119.237e-18
c2982 n176__vddio vss 101.022e-18
c2983 n177__vddio vss 129.788e-18
c2984 n178__vddio vss 98.228e-18
c2985 n1161__vddio vss 54.6006e-18
c2986 n170__i1__i14__net1 vss 39.4314e-18
c2987 n6__i5__i7__x0out vss 70.6656e-18
c2988 n299__chipdriverout vss 101.362e-18
c2989 n300__chipdriverout vss 121.262e-18
c2990 n301__chipdriverout vss 121.085e-18
c2991 n302__chipdriverout vss 105.597e-18
c2992 n303__chipdriverout vss 89.6537e-18
c2993 n304__chipdriverout vss 92.2442e-18
c2994 n305__chipdriverout vss 104.17e-18
c2995 n306__chipdriverout vss 119.104e-18
c2996 n307__chipdriverout vss 120.275e-18
c2997 n308__chipdriverout vss 107.347e-18
c2998 n309__chipdriverout vss 125.955e-18
c2999 n310__chipdriverout vss 124.268e-18
c3000 n311__chipdriverout vss 124.234e-18
c3001 n167__i1__i14__net1 vss 40.615e-18
c3002 n11__reset vss 24.0848e-18
c3003 n10__reset vss 22.5356e-18
c3004 n151__vddio vss 121.331e-18
c3005 n152__vddio vss 119.408e-18
c3006 n153__vddio vss 120.253e-18
c3007 n154__vddio vss 119.323e-18
c3008 n155__vddio vss 117.031e-18
c3009 n156__vddio vss 113.436e-18
c3010 n157__vddio vss 113.038e-18
c3011 n1162__vddio vss 75.5506e-18
c3012 n155__i1__i14__net1 vss 39.3708e-18
c3013 n260__chipdriverout vss 101.498e-18
c3014 n261__chipdriverout vss 121.262e-18
c3015 n262__chipdriverout vss 137.457e-18
c3016 n263__chipdriverout vss 121.738e-18
c3017 n264__chipdriverout vss 89.6537e-18
c3018 n265__chipdriverout vss 92.2612e-18
c3019 n266__chipdriverout vss 120.096e-18
c3020 n267__chipdriverout vss 135.498e-18
c3021 n268__chipdriverout vss 120.304e-18
c3022 n269__chipdriverout vss 106.301e-18
c3023 n270__chipdriverout vss 124.39e-18
c3024 n271__chipdriverout vss 122.347e-18
c3025 n272__chipdriverout vss 126.311e-18
c3026 n151__i1__i14__net1 vss 40.7527e-18
c3027 n66__vdd vss 103.34e-18
c3028 n130__vddio vss 121.42e-18
c3029 n131__vddio vss 119.588e-18
c3030 n132__vddio vss 120.348e-18
c3031 n133__vddio vss 119.431e-18
c3032 n134__vddio vss 117.128e-18
c3033 n135__vddio vss 114.714e-18
c3034 n136__vddio vss 115.031e-18
c3035 n1163__vddio vss 54.7056e-18
c3036 n139__i1__i14__net1 vss 40.9087e-18
c3037 n221__chipdriverout vss 102.307e-18
c3038 n222__chipdriverout vss 122.701e-18
c3039 n223__chipdriverout vss 139.11e-18
c3040 n224__chipdriverout vss 123.186e-18
c3041 n225__chipdriverout vss 90.5284e-18
c3042 n226__chipdriverout vss 92.622e-18
c3043 n227__chipdriverout vss 122.102e-18
c3044 n228__chipdriverout vss 137.875e-18
c3045 n229__chipdriverout vss 122.316e-18
c3046 n230__chipdriverout vss 107.541e-18
c3047 n231__chipdriverout vss 124.975e-18
c3048 n232__chipdriverout vss 122.207e-18
c3049 n233__chipdriverout vss 130.099e-18
c3050 n135__i1__i14__net1 vss 39.743e-18
c3051 n109__vddio vss 120.913e-18
c3052 n110__vddio vss 118.829e-18
c3053 n111__vddio vss 119.841e-18
c3054 n112__vddio vss 118.955e-18
c3055 n113__vddio vss 116.674e-18
c3056 n114__vddio vss 114.005e-18
c3057 n115__vddio vss 114.578e-18
c3058 n1164__vddio vss 77.4007e-18
c3059 n15__i5__i7__i1__net1 vss 154.837e-18
c3060 n15__i5__i7__i0__net1 vss 287.594e-18
c3061 n121__i1__i14__net1 vss 40.8198e-18
c3062 n182__chipdriverout vss 101.041e-18
c3063 n183__chipdriverout vss 120.679e-18
c3064 n184__chipdriverout vss 137.002e-18
c3065 n185__chipdriverout vss 121.152e-18
c3066 n186__chipdriverout vss 89.323e-18
c3067 n187__chipdriverout vss 91.279e-18
c3068 n188__chipdriverout vss 119.683e-18
c3069 n189__chipdriverout vss 135.148e-18
c3070 n190__chipdriverout vss 119.889e-18
c3071 n191__chipdriverout vss 105.096e-18
c3072 n192__chipdriverout vss 122.488e-18
c3073 n193__chipdriverout vss 119.457e-18
c3074 n194__chipdriverout vss 127.759e-18
c3075 n1595__vddio vss 11.1885e-18
c3076 n119__i1__i14__net1 vss 42.4887e-18
c3077 n7__y0 vss 15.4912e-18
c3078 n7__x0 vss 13.2076e-18
c3079 n82__vddio vss 103.564e-18
c3080 n83__vddio vss 135.767e-18
c3081 n84__vddio vss 104.339e-18
c3082 n85__vddio vss 103.163e-18
c3083 n86__vddio vss 100.913e-18
c3084 n87__vddio vss 130.893e-18
c3085 n88__vddio vss 99.0364e-18
c3086 n1165__vddio vss 54.2498e-18
c3087 n111__i1__i14__net1 vss 39.7359e-18
c3088 n143__chipdriverout vss 116.272e-18
c3089 n144__chipdriverout vss 103.26e-18
c3090 n145__chipdriverout vss 118.883e-18
c3091 n146__chipdriverout vss 103.525e-18
c3092 n147__chipdriverout vss 69.6341e-18
c3093 n148__chipdriverout vss 112.584e-18
c3094 n149__chipdriverout vss 102.452e-18
c3095 n150__chipdriverout vss 117.21e-18
c3096 n151__chipdriverout vss 102.452e-18
c3097 n152__chipdriverout vss 119.784e-18
c3098 n153__chipdriverout vss 105.22e-18
c3099 n154__chipdriverout vss 134.083e-18
c3100 n155__chipdriverout vss 109.783e-18
c3101 n10__i5__i7__i1__net1 vss 96.4527e-18
c3102 n10__i5__i7__i0__net1 vss 93.0607e-18
c3103 n103__i1__i14__net1 vss 40.7164e-18
c3104 n57__vddio vss 103.799e-18
c3105 n58__vddio vss 135.649e-18
c3106 n59__vddio vss 104.445e-18
c3107 n60__vddio vss 103.274e-18
c3108 n61__vddio vss 101.02e-18
c3109 n62__vddio vss 130.774e-18
c3110 n63__vddio vss 99.1422e-18
c3111 n1166__vddio vss 54.5737e-18
c3112 n95__i1__i14__net1 vss 41.3494e-18
c3113 n19__i5__clk4 vss 100.325e-18
c3114 n104__chipdriverout vss 142.68e-18
c3115 n105__chipdriverout vss 108.096e-18
c3116 n106__chipdriverout vss 121.593e-18
c3117 n107__chipdriverout vss 109.035e-18
c3118 n108__chipdriverout vss 71.3167e-18
c3119 n109__chipdriverout vss 114.612e-18
c3120 n110__chipdriverout vss 104.435e-18
c3121 n111__chipdriverout vss 119.398e-18
c3122 n112__chipdriverout vss 104.435e-18
c3123 n113__chipdriverout vss 121.829e-18
c3124 n114__chipdriverout vss 107.659e-18
c3125 n115__chipdriverout vss 136.353e-18
c3126 n116__chipdriverout vss 111.694e-18
c3127 n85__i1__i14__net1 vss 42.6763e-18
c3128 n36__vddio vss 103.764e-18
c3129 n37__vddio vss 135.649e-18
c3130 n38__vddio vss 104.445e-18
c3131 n39__vddio vss 103.274e-18
c3132 n40__vddio vss 101.02e-18
c3133 n41__vddio vss 129.83e-18
c3134 n42__vddio vss 98.225e-18
c3135 n1167__vddio vss 76.357e-18
c3136 n75__i1__i14__net1 vss 40.4563e-18
c3137 n65__chipdriverout vss 136.955e-18
c3138 n66__chipdriverout vss 110.156e-18
c3139 n67__chipdriverout vss 127.342e-18
c3140 n68__chipdriverout vss 110.405e-18
c3141 n69__chipdriverout vss 73.5898e-18
c3142 n70__chipdriverout vss 116.57e-18
c3143 n71__chipdriverout vss 106.66e-18
c3144 n72__chipdriverout vss 119.398e-18
c3145 n73__chipdriverout vss 104.435e-18
c3146 n74__chipdriverout vss 126.487e-18
c3147 n75__chipdriverout vss 109.785e-18
c3148 n76__chipdriverout vss 141.737e-18
c3149 n77__chipdriverout vss 107.215e-18
c3150 n71__i1__i14__net1 vss 43.1823e-18
c3151 n15__vddio vss 72.7535e-18
c3152 n16__vddio vss 104.859e-18
c3153 n17__vddio vss 73.4856e-18
c3154 n18__vddio vss 75.4059e-18
c3155 n19__vddio vss 76.5607e-18
c3156 n20__vddio vss 106.465e-18
c3157 n21__vddio vss 74.175e-18
c3158 n63__i1__i14__net1 vss 70.6503e-18
c3159 n26__chipdriverout vss 57.1757e-18
c3160 n27__chipdriverout vss 39.2247e-18
c3161 n28__chipdriverout vss 40.3569e-18
c3162 n29__chipdriverout vss 40.0826e-18
c3163 n30__chipdriverout vss 34.2978e-18
c3164 n31__chipdriverout vss 60.6769e-18
c3165 n32__chipdriverout vss 34.5734e-18
c3166 n33__chipdriverout vss 40.6968e-18
c3167 n34__chipdriverout vss 37.5967e-18
c3168 n35__chipdriverout vss 44.0422e-18
c3169 n36__chipdriverout vss 40.424e-18
c3170 n37__chipdriverout vss 51.8943e-18
c3171 n38__chipdriverout vss 49.2191e-18
c3172 n1819__vddio vss 129.397e-18
c3173 n1817__vddio vss 150.715e-18
c3174 n1814__vddio vss 101.934e-18
c3175 n1820__vddio vss 3.81878e-18
c3176 n1813__vddio vss 69.6313e-18
c3177 n64__i1__net3 vss 60.972e-18
c3178 n65__i1__net3 vss 44.8286e-18
c3179 n182__i1__i13__net1 vss 268.524e-18
c3180 n184__i1__i13__net1 vss 328.873e-18
c3181 n190__i1__i13__net1 vss 237.381e-18
c3182 n189__i1__i13__net1 vss 276.629e-18
c3183 n186__i1__i13__net1 vss 296.549e-18
c3184 n62__i1__net3 vss 61.1232e-18
c3185 n63__i1__net3 vss 40.6013e-18
c3186 n1806__vddio vss 256.815e-18
c3187 n1809__vddio vss 342.389e-18
c3188 n1811__vddio vss 251.259e-18
c3189 n1812__vddio vss 152.923e-18
c3190 n60__i1__net3 vss 61.1267e-18
c3191 n61__i1__net3 vss 38.8384e-18
c3192 n171__i1__i13__net1 vss 281.779e-18
c3193 n173__i1__i13__net1 vss 347.149e-18
c3194 n179__i1__i13__net1 vss 258.074e-18
c3195 n178__i1__i13__net1 vss 297.303e-18
c3196 n175__i1__i13__net1 vss 329.398e-18
c3197 n58__i1__net3 vss 61.2688e-18
c3198 n59__i1__net3 vss 40.7254e-18
c3199 n1799__vddio vss 264.724e-18
c3200 n1802__vddio vss 345.084e-18
c3201 n1804__vddio vss 252.342e-18
c3202 n1805__vddio vss 152.205e-18
c3203 n56__i1__net3 vss 61.5786e-18
c3204 n57__i1__net3 vss 39.7944e-18
c3205 n160__i1__i13__net1 vss 280.81e-18
c3206 n162__i1__i13__net1 vss 341.705e-18
c3207 n168__i1__i13__net1 vss 257.867e-18
c3208 n167__i1__i13__net1 vss 295.314e-18
c3209 n164__i1__i13__net1 vss 314.09e-18
c3210 n54__i1__net3 vss 74.6078e-18
c3211 n55__i1__net3 vss 48.283e-18
c3212 n1798__vddio vss 198.325e-18
c3213 n1796__vddio vss 287.782e-18
c3214 n1793__vddio vss 226.504e-18
c3215 n1792__vddio vss 123.065e-18
c3216 n1822__vddio vss 3.56162e-18
c3217 n1785__vddio vss 169.119e-18
c3218 n1788__vddio vss 192.839e-18
c3219 n1790__vddio vss 144.831e-18
c3220 n1791__vddio vss 85.4602e-18
c3221 n157__i1__i13__net1 vss 43.4095e-18
c3222 n158__i1__i13__net1 vss 37.9704e-18
c3223 n324__i1__net2 vss 275.65e-18
c3224 n325__i1__net2 vss 278.59e-18
c3225 n328__i1__net2 vss 308.684e-18
c3226 n17__piso_outinv vss 90.4464e-18
c3227 n11__i1__i11__outinv vss 306.298e-18
c3228 n321__i1__net2 vss 266.574e-18
c3229 n323__i1__net2 vss 312.399e-18
c3230 n25__i1__net4 vss 275.904e-18
c3231 n155__i1__i13__net1 vss 64.149e-18
c3232 n156__i1__i13__net1 vss 52.9451e-18
c3233 n16__piso_outinv vss 59.1041e-18
c3234 n1759__vddio vss 265.137e-18
c3235 n1762__vddio vss 347.572e-18
c3236 n1764__vddio vss 250.387e-18
c3237 n1765__vddio vss 156.423e-18
c3238 n10__i1__i11__outinv vss 105.663e-18
c3239 n153__i1__i13__net1 vss 54.2808e-18
c3240 n154__i1__i13__net1 vss 34.9382e-18
c3241 n315__i1__net2 vss 293.892e-18
c3242 n316__i1__net2 vss 297.877e-18
c3243 n319__i1__net2 vss 327.984e-18
c3244 n15__piso_outinv vss 111.735e-18
c3245 n312__i1__net2 vss 291.507e-18
c3246 n314__i1__net2 vss 339.147e-18
c3247 n151__i1__i13__net1 vss 64.242e-18
c3248 n152__i1__i13__net1 vss 36.0103e-18
c3249 n1752__vddio vss 268.603e-18
c3250 n1755__vddio vss 349.391e-18
c3251 n1757__vddio vss 253.168e-18
c3252 n1758__vddio vss 151.662e-18
c3253 n149__i1__i13__net1 vss 31.9778e-18
c3254 n150__i1__i13__net1 vss 53.0975e-18
c3255 n308__i1__net2 vss 290.786e-18
c3256 n310__i1__net2 vss 339.985e-18
c3257 n302__i1__net2 vss 316.591e-18
c3258 n303__i1__net2 vss 303.766e-18
c3259 n306__i1__net2 vss 333.709e-18
c3260 n23__i1__net4 vss 69.8587e-18
c3261 n1745__vddio vss 268.65e-18
c3262 n1748__vddio vss 352.044e-18
c3263 n1750__vddio vss 254.541e-18
c3264 n1751__vddio vss 114.627e-18
c3265 n31__piso_out vss 84.957e-18
c3266 n141__i1__i13__net1 vss 64.4841e-18
c3267 n142__i1__i13__net1 vss 53.1317e-18
c3268 n299__i1__net2 vss 290.001e-18
c3269 n301__i1__net2 vss 347.113e-18
c3270 n293__i1__net2 vss 296.839e-18
c3271 n294__i1__net2 vss 300.667e-18
c3272 n297__i1__net2 vss 332.561e-18
c3273 n22__i1__net4 vss 93.6195e-18
c3274 n28__piso_out vss 82.7112e-18
c3275 n137__i1__i13__net1 vss 63.7365e-18
c3276 n138__i1__i13__net1 vss 35.9854e-18
c3277 n7__i1__i11__outinv vss 268.866e-18
c3278 n1738__vddio vss 265.539e-18
c3279 n1741__vddio vss 350.844e-18
c3280 n1743__vddio vss 257.102e-18
c3281 n1744__vddio vss 155.071e-18
c3282 n133__i1__i13__net1 vss 41.4617e-18
c3283 n134__i1__i13__net1 vss 52.0809e-18
c3284 n1730__vddio vss 26.6648e-18
c3285 n290__i1__net2 vss 285.487e-18
c3286 n292__i1__net2 vss 344.39e-18
c3287 n284__i1__net2 vss 292.17e-18
c3288 n285__i1__net2 vss 295.01e-18
c3289 n288__i1__net2 vss 328.148e-18
c3290 n129__i1__i13__net1 vss 41.0845e-18
c3291 n130__i1__i13__net1 vss 53.0088e-18
c3292 n17__i1__net4 vss 46.5763e-18
c3293 n18__i1__net4 vss 44.7353e-18
c3294 n1713__vddio vss 266.752e-18
c3295 n1716__vddio vss 348.755e-18
c3296 n1718__vddio vss 252.89e-18
c3297 n1719__vddio vss 153.321e-18
c3298 n125__i1__i13__net1 vss 64.3666e-18
c3299 n126__i1__i13__net1 vss 52.0809e-18
c3300 n65__i1__i12__net1 vss 319.243e-18
c3301 n64__i1__i12__net1 vss 266.045e-18
c3302 n281__i1__net2 vss 284.72e-18
c3303 n283__i1__net2 vss 344.655e-18
c3304 n275__i1__net2 vss 292.661e-18
c3305 n276__i1__net2 vss 298.498e-18
c3306 n279__i1__net2 vss 333.369e-18
c3307 n13__i1__net4 vss 78.6709e-18
c3308 n14__i1__net4 vss 46.5547e-18
c3309 n117__i1__i13__net1 vss 40.7445e-18
c3310 n118__i1__i13__net1 vss 53.1099e-18
c3311 n1712__vddio vss 268.955e-18
c3312 n1710__vddio vss 348.149e-18
c3313 n1707__vddio vss 248.862e-18
c3314 n1706__vddio vss 168e-18
c3315 n113__i1__i13__net1 vss 40.2372e-18
c3316 n114__i1__i13__net1 vss 54.6407e-18
c3317 n1733__vddio vss 34.9402e-18
c3318 n272__i1__net2 vss 301.192e-18
c3319 n274__i1__net2 vss 355.623e-18
c3320 n266__i1__net2 vss 313.512e-18
c3321 n267__i1__net2 vss 312.369e-18
c3322 n270__i1__net2 vss 336.103e-18
c3323 n1826__vddio vss 83.346e-18
c3324 n1699__vddio vss 254.243e-18
c3325 n1702__vddio vss 343.249e-18
c3326 n1704__vddio vss 248.759e-18
c3327 n1705__vddio vss 153.369e-18
c3328 n28__i1__net3 vss 76.7887e-18
c3329 n26__i1__net3 vss 225.457e-18
c3330 n263__i1__net2 vss 284.858e-18
c3331 n265__i1__net2 vss 339.037e-18
c3332 n257__i1__net2 vss 293.952e-18
c3333 n258__i1__net2 vss 297.828e-18
c3334 n261__i1__net2 vss 325.361e-18
c3335 n49__i1__i12__net1 vss 35.0372e-18
c3336 n50__i1__i12__net1 vss 46.8754e-18
c3337 n101__i1__i13__net1 vss 41.0286e-18
c3338 n102__i1__i13__net1 vss 52.9383e-18
c3339 n1692__vddio vss 252.626e-18
c3340 n1695__vddio vss 339.666e-18
c3341 n1697__vddio vss 244.194e-18
c3342 n1698__vddio vss 152.218e-18
c3343 n45__i1__i12__net1 vss 54.9991e-18
c3344 n46__i1__i12__net1 vss 31.6537e-18
c3345 n21__i1__net3 vss 237.876e-18
c3346 n17__i1__net3 vss 270.443e-18
c3347 n254__i1__net2 vss 285.778e-18
c3348 n256__i1__net2 vss 339.373e-18
c3349 n248__i1__net2 vss 296.449e-18
c3350 n249__i1__net2 vss 300.073e-18
c3351 n252__i1__net2 vss 326.594e-18
c3352 n41__i1__i12__net1 vss 58.5643e-18
c3353 n42__i1__i12__net1 vss 34.5034e-18
c3354 n85__i1__i13__net1 vss 63.4774e-18
c3355 n86__i1__i13__net1 vss 36.6623e-18
c3356 n1685__vddio vss 261.721e-18
c3357 n1688__vddio vss 348.875e-18
c3358 n1690__vddio vss 251.672e-18
c3359 n1691__vddio vss 153.125e-18
c3360 n37__i1__i12__net1 vss 58.8819e-18
c3361 n38__i1__i12__net1 vss 37.3467e-18
c3362 n73__i1__i13__net1 vss 63.3152e-18
c3363 n74__i1__i13__net1 vss 34.984e-18
c3364 n8__i1__net3 vss 283.971e-18
c3365 n14__i1__net3 vss 242.981e-18
c3366 n243__i1__net2 vss 309.167e-18
c3367 n244__i1__net2 vss 304.848e-18
c3368 n247__i1__net2 vss 333.347e-18
c3369 n240__i1__net2 vss 300.269e-18
c3370 n242__i1__net2 vss 357.971e-18
c3371 n33__i1__i12__net1 vss 35.7497e-18
c3372 n34__i1__i12__net1 vss 41.177e-18
c3373 n1678__vddio vss 254.897e-18
c3374 n1681__vddio vss 333.973e-18
c3375 n1683__vddio vss 242.96e-18
c3376 n1684__vddio vss 139.122e-18
c3377 n29__i1__i12__net1 vss 47.8658e-18
c3378 n30__i1__i12__net1 vss 69.9871e-18
c3379 n61__i1__i13__net1 vss 51.6584e-18
c3380 n62__i1__i13__net1 vss 63.1698e-18
c3381 n6__i1__net3 vss 139.299e-18
c3382 n236__i1__net2 vss 140.741e-18
c3383 n238__i1__net2 vss 173.923e-18
c3384 n230__i1__net2 vss 134.005e-18
c3385 n231__i1__net2 vss 139.152e-18
c3386 n234__i1__net2 vss 185.699e-18
c3387 n184__vdd vss 74.4012e-18
c3388 n1494__vddio vss 163.419e-18
c3389 n1495__vddio vss 153.31e-18
c3390 n1498__vddio vss 80.6754e-18
c3391 n1499__vddio vss 154.175e-18
c3392 n1502__vddio vss 80.8779e-18
c3393 n1503__vddio vss 148.813e-18
c3394 n1506__vddio vss 80.0447e-18
c3395 n221__i1__net2 vss 44.8678e-18
c3396 n222__i1__net2 vss 54.7533e-18
c3397 n45__shift vss 63.7218e-18
c3398 n1298__i1__i14__net1 vss 131.363e-18
c3399 n1301__i1__i14__net1 vss 226.368e-18
c3400 n1302__i1__i14__net1 vss 195.211e-18
c3401 n1305__i1__i14__net1 vss 232.194e-18
c3402 n1306__i1__i14__net1 vss 273.678e-18
c3403 n1309__i1__i14__net1 vss 228.936e-18
c3404 n1310__i1__i14__net1 vss 200.135e-18
c3405 n1313__i1__i14__net1 vss 226.434e-18
c3406 n1314__i1__i14__net1 vss 204.434e-18
c3407 n1317__i1__i14__net1 vss 202.713e-18
c3408 n1318__i1__i14__net1 vss 198.275e-18
c3409 n1321__i1__i14__net1 vss 203.721e-18
c3410 n1322__i1__i14__net1 vss 254.196e-18
c3411 n217__i1__net2 vss 43.4541e-18
c3412 n218__i1__net2 vss 37.0267e-18
c3413 n2__piso_outinv vss 57.9802e-18
c3414 n1473__vddio vss 272.092e-18
c3415 n1474__vddio vss 257.805e-18
c3416 n1477__vddio vss 136.37e-18
c3417 n1478__vddio vss 245.986e-18
c3418 n1481__vddio vss 141.624e-18
c3419 n1482__vddio vss 256.353e-18
c3420 n1485__vddio vss 140.285e-18
c3421 n1492__vddio vss 164.878e-18
c3422 n1262__i1__i14__net1 vss 144.986e-18
c3423 n1263__i1__i14__net1 vss 203.238e-18
c3424 n1265__i1__i14__net1 vss 171.36e-18
c3425 n1266__i1__i14__net1 vss 208.697e-18
c3426 n1268__i1__i14__net1 vss 247.008e-18
c3427 n1271__i1__i14__net1 vss 253.613e-18
c3428 n1274__i1__i14__net1 vss 177.144e-18
c3429 n1275__i1__i14__net1 vss 200.637e-18
c3430 n1277__i1__i14__net1 vss 178.932e-18
c3431 n1278__i1__i14__net1 vss 220.105e-18
c3432 n1280__i1__i14__net1 vss 173.382e-18
c3433 n1281__i1__i14__net1 vss 220.562e-18
c3434 n1283__i1__i14__net1 vss 229.23e-18
c3435 n37__i5__i8__net2 vss 68.1795e-18
c3436 n209__i1__net2 vss 36.3503e-18
c3437 n210__i1__net2 vss 47.9251e-18
c3438 n101__i5__clk4 vss 88.1358e-18
c3439 n1533__vddio vss 5.31338e-18
c3440 n1452__vddio vss 284.401e-18
c3441 n1455__vddio vss 237.523e-18
c3442 n1456__vddio vss 150.988e-18
c3443 n1458__vddio vss 258.132e-18
c3444 n1459__vddio vss 156.159e-18
c3445 n1461__vddio vss 236.718e-18
c3446 n1462__vddio vss 154.986e-18
c3447 n1464__vddio vss 187.296e-18
c3448 n205__i1__net2 vss 39.1038e-18
c3449 n206__i1__net2 vss 47.7041e-18
c3450 n1238__i1__i14__net1 vss 143.357e-18
c3451 n1239__i1__i14__net1 vss 201.365e-18
c3452 n1241__i1__i14__net1 vss 171.05e-18
c3453 n1242__i1__i14__net1 vss 206.422e-18
c3454 n1244__i1__i14__net1 vss 246.9e-18
c3455 n1221__i1__i14__net1 vss 256.97e-18
c3456 n1224__i1__i14__net1 vss 183.389e-18
c3457 n1225__i1__i14__net1 vss 208.869e-18
c3458 n1227__i1__i14__net1 vss 185.315e-18
c3459 n1228__i1__i14__net1 vss 228.279e-18
c3460 n1230__i1__i14__net1 vss 179.29e-18
c3461 n1231__i1__i14__net1 vss 228.678e-18
c3462 n1233__i1__i14__net1 vss 233.327e-18
c3463 n11__i5__i8__net5 vss 54.7661e-18
c3464 n201__i1__net2 vss 36.3503e-18
c3465 n202__i1__net2 vss 46.4967e-18
c3466 n1431__vddio vss 264.406e-18
c3467 n1434__vddio vss 251.819e-18
c3468 n1435__vddio vss 133.724e-18
c3469 n1437__vddio vss 239.632e-18
c3470 n1438__vddio vss 138.706e-18
c3471 n1440__vddio vss 250.972e-18
c3472 n1441__vddio vss 137.686e-18
c3473 n1443__vddio vss 161.851e-18
c3474 n197__i1__net2 vss 46.2309e-18
c3475 n198__i1__net2 vss 38.6665e-18
c3476 n1199__i1__i14__net1 vss 128.033e-18
c3477 n1200__i1__i14__net1 vss 218.316e-18
c3478 n1202__i1__i14__net1 vss 187.504e-18
c3479 n1203__i1__i14__net1 vss 224.256e-18
c3480 n1205__i1__i14__net1 vss 265.466e-18
c3481 n1182__i1__i14__net1 vss 231.09e-18
c3482 n1185__i1__i14__net1 vss 196.565e-18
c3483 n1186__i1__i14__net1 vss 222.476e-18
c3484 n1188__i1__i14__net1 vss 198.782e-18
c3485 n1189__i1__i14__net1 vss 209.447e-18
c3486 n1191__i1__i14__net1 vss 192.513e-18
c3487 n1192__i1__i14__net1 vss 209.827e-18
c3488 n1194__i1__i14__net1 vss 249.305e-18
c3489 n193__i1__net2 vss 36.3332e-18
c3490 n194__i1__net2 vss 35.6393e-18
c3491 n94__i5__clk4 vss 49.5587e-18
c3492 n1410__vddio vss 288.578e-18
c3493 n1413__vddio vss 238.698e-18
c3494 n1414__vddio vss 150.503e-18
c3495 n1416__vddio vss 259.017e-18
c3496 n1417__vddio vss 155.93e-18
c3497 n1419__vddio vss 237.206e-18
c3498 n1420__vddio vss 154.348e-18
c3499 n1422__vddio vss 184.707e-18
c3500 n189__i1__net2 vss 46.1183e-18
c3501 n190__i1__net2 vss 39.7462e-18
c3502 n1145__i1__i14__net1 vss 16.1516e-18
c3503 n1146__i1__i14__net1 vss 202.357e-18
c3504 n1148__i1__i14__net1 vss 171.251e-18
c3505 n1149__i1__i14__net1 vss 208.208e-18
c3506 n1151__i1__i14__net1 vss 246.909e-18
c3507 n1154__i1__i14__net1 vss 250.334e-18
c3508 n1157__i1__i14__net1 vss 174.603e-18
c3509 n1158__i1__i14__net1 vss 197.995e-18
c3510 n1160__i1__i14__net1 vss 176.481e-18
c3511 n1161__i1__i14__net1 vss 217.193e-18
c3512 n1163__i1__i14__net1 vss 170.804e-18
c3513 n1164__i1__i14__net1 vss 218.049e-18
c3514 n1166__i1__i14__net1 vss 226.601e-18
c3515 n1379__vddio vss 274.949e-18
c3516 n1382__vddio vss 240.709e-18
c3517 n1383__vddio vss 135.969e-18
c3518 n1385__vddio vss 245.191e-18
c3519 n1386__vddio vss 157.218e-18
c3520 n1388__vddio vss 239.016e-18
c3521 n1389__vddio vss 154.391e-18
c3522 n1391__vddio vss 163.263e-18
c3523 n69__reset vss 59.5418e-18
c3524 n68__reset vss 85.1574e-18
c3525 n177__i1__net2 vss 39.0801e-18
c3526 n178__i1__net2 vss 48.9234e-18
c3527 n9__i5__i8__i10__net24 vss 62.4343e-18
c3528 n6__i5__i8__i10__net23 vss 84.833e-18
c3529 n7__i5__i6__i5__net24 vss 50.6624e-18
c3530 n6__i5__i6__i5__net23 vss 77.5023e-18
c3531 n1106__i1__i14__net1 vss 128.055e-18
c3532 n1107__i1__i14__net1 vss 218.194e-18
c3533 n1109__i1__i14__net1 vss 187.504e-18
c3534 n1110__i1__i14__net1 vss 224.256e-18
c3535 n1112__i1__i14__net1 vss 265.473e-18
c3536 n1115__i1__i14__net1 vss 230.604e-18
c3537 n1118__i1__i14__net1 vss 193.014e-18
c3538 n1119__i1__i14__net1 vss 216.945e-18
c3539 n1121__i1__i14__net1 vss 195.008e-18
c3540 n1122__i1__i14__net1 vss 203.995e-18
c3541 n1124__i1__i14__net1 vss 188.944e-18
c3542 n1125__i1__i14__net1 vss 203.723e-18
c3543 n1127__i1__i14__net1 vss 245.016e-18
c3544 n171__i1__net2 vss 23.7365e-18
c3545 n172__i1__net2 vss 48.0997e-18
c3546 n27__i5__i8__net1 vss 260.211e-18
c3547 n35__i5__i8__net2 vss 122.798e-18
c3548 n44__i5__i6__net31 vss 227.24e-18
c3549 n67__i5__clk_buf vss 120.425e-18
c3550 n6__i5__i8__i10__net24 vss 109.123e-18
c3551 n3__i5__i8__i10__net23 vss 97.3471e-18
c3552 n1358__vddio vss 266.24e-18
c3553 n1361__vddio vss 253.929e-18
c3554 n1362__vddio vss 135.016e-18
c3555 n1364__vddio vss 241.917e-18
c3556 n1365__vddio vss 139.984e-18
c3557 n1367__vddio vss 252.956e-18
c3558 n1368__vddio vss 138.743e-18
c3559 n1370__vddio vss 164.455e-18
c3560 n6__i5__i6__i5__net24 vss 105.523e-18
c3561 n3__i5__i6__i5__net23 vss 98.4925e-18
c3562 n169__i1__net2 vss 46.1359e-18
c3563 n170__i1__net2 vss 38.6298e-18
c3564 n1064__i1__i14__net1 vss 128.033e-18
c3565 n1067__i1__i14__net1 vss 218.194e-18
c3566 n1068__i1__i14__net1 vss 187.504e-18
c3567 n1071__i1__i14__net1 vss 224.256e-18
c3568 n1072__i1__i14__net1 vss 265.473e-18
c3569 n1075__i1__i14__net1 vss 234.244e-18
c3570 n1076__i1__i14__net1 vss 199.196e-18
c3571 n1079__i1__i14__net1 vss 225.115e-18
c3572 n1080__i1__i14__net1 vss 201.33e-18
c3573 n1083__i1__i14__net1 vss 212.229e-18
c3574 n1084__i1__i14__net1 vss 195.097e-18
c3575 n1087__i1__i14__net1 vss 212.431e-18
c3576 n1088__i1__i14__net1 vss 251.143e-18
c3577 n3__i5__i8__i10__net24 vss 106.723e-18
c3578 n2__i5__i8__i10__net23 vss 107.444e-18
c3579 n3__i5__i6__i5__net24 vss 103.459e-18
c3580 n2__i5__i6__i5__net23 vss 106.562e-18
c3581 n1336__vddio vss 281.7e-18
c3582 n1339__vddio vss 235.452e-18
c3583 n1340__vddio vss 149.598e-18
c3584 n1343__vddio vss 255.747e-18
c3585 n1344__vddio vss 154.782e-18
c3586 n1347__vddio vss 234.605e-18
c3587 n1348__vddio vss 153.543e-18
c3588 n1356__vddio vss 185.119e-18
c3589 n7__i5__i8__i10__net25 vss 102.74e-18
c3590 n6__i5__i8__i10__net21 vss 110.07e-18
c3591 n7__i5__i6__i5__net25 vss 103.224e-18
c3592 n6__i5__i6__i5__net21 vss 107.004e-18
c3593 n1043__i1__i14__net1 vss 134.257e-18
c3594 n1044__i1__i14__net1 vss 223.962e-18
c3595 n1046__i1__i14__net1 vss 176.602e-18
c3596 n1047__i1__i14__net1 vss 229.458e-18
c3597 n1049__i1__i14__net1 vss 269.317e-18
c3598 n1026__i1__i14__net1 vss 235.159e-18
c3599 n1029__i1__i14__net1 vss 201.32e-18
c3600 n1030__i1__i14__net1 vss 228.38e-18
c3601 n1032__i1__i14__net1 vss 203.714e-18
c3602 n1033__i1__i14__net1 vss 215.252e-18
c3603 n1035__i1__i14__net1 vss 197.221e-18
c3604 n1036__i1__i14__net1 vss 215.931e-18
c3605 n1038__i1__i14__net1 vss 256.492e-18
c3606 n26__i5__i8__net1 vss 286.798e-18
c3607 n33__i5__i8__net2 vss 363.822e-18
c3608 n41__i5__i6__net31 vss 118.497e-18
c3609 n65__i5__clk_buf vss 144.555e-18
c3610 n6__i5__i8__i10__net25 vss 116.396e-18
c3611 n3__i5__i8__i10__net21 vss 91.3919e-18
c3612 n6__i5__i6__i5__net25 vss 115.912e-18
c3613 n3__i5__i6__i5__net21 vss 88.3067e-18
c3614 n157__i1__net2 vss 45.1816e-18
c3615 n158__i1__net2 vss 37.296e-18
c3616 n194__vdd vss 104.819e-18
c3617 n8__i5__i8__net5 vss 32.6165e-18
c3618 n1316__vddio vss 267.229e-18
c3619 n1319__vddio vss 254.279e-18
c3620 n1320__vddio vss 134.175e-18
c3621 n1322__vddio vss 241.835e-18
c3622 n1323__vddio vss 139.565e-18
c3623 n1325__vddio vss 253.377e-18
c3624 n1326__vddio vss 137.995e-18
c3625 n1328__vddio vss 184.572e-18
c3626 n3__i5__i8__i10__net25 vss 89.2432e-18
c3627 n2__i5__i8__i10__net21 vss 114.041e-18
c3628 n149__i1__net2 vss 46.4869e-18
c3629 n150__i1__net2 vss 39.1206e-18
c3630 n3__i5__i6__i5__net25 vss 82.5929e-18
c3631 n2__i5__i6__i5__net21 vss 93.4228e-18
c3632 n15__i5__i6__net35 vss 69.4921e-18
c3633 n989__i1__i14__net1 vss 135.089e-18
c3634 n990__i1__i14__net1 vss 228.68e-18
c3635 n992__i1__i14__net1 vss 196.575e-18
c3636 n993__i1__i14__net1 vss 234.038e-18
c3637 n995__i1__i14__net1 vss 274.311e-18
c3638 n998__i1__i14__net1 vss 230.267e-18
c3639 n1001__i1__i14__net1 vss 194.603e-18
c3640 n1002__i1__i14__net1 vss 218.535e-18
c3641 n1004__i1__i14__net1 vss 196.612e-18
c3642 n1005__i1__i14__net1 vss 205.482e-18
c3643 n1007__i1__i14__net1 vss 190.842e-18
c3644 n1008__i1__i14__net1 vss 205.731e-18
c3645 n1010__i1__i14__net1 vss 246.467e-18
c3646 n19__i5__i8__net1 vss 122.231e-18
c3647 n141__i1__net2 vss 35.737e-18
c3648 n142__i1__net2 vss 47.5703e-18
c3649 n9__i5__i6__net35 vss 59.0223e-18
c3650 n1295__vddio vss 288.409e-18
c3651 n1298__vddio vss 240.65e-18
c3652 n1299__vddio vss 151.776e-18
c3653 n1301__vddio vss 261.211e-18
c3654 n1302__vddio vss 157.187e-18
c3655 n1304__vddio vss 239.198e-18
c3656 n1305__vddio vss 155.673e-18
c3657 n1307__vddio vss 164.34e-18
c3658 n12__i5__r0 vss 96.2133e-18
c3659 n129__i1__net2 vss 39.2353e-18
c3660 n130__i1__net2 vss 47.043e-18
c3661 n951__i1__i14__net1 vss 229.9e-18
c3662 n953__i1__i14__net1 vss 196.891e-18
c3663 n954__i1__i14__net1 vss 236.094e-18
c3664 n956__i1__i14__net1 vss 274.512e-18
c3665 n959__i1__i14__net1 vss 226.039e-18
c3666 n962__i1__i14__net1 vss 190.993e-18
c3667 n963__i1__i14__net1 vss 214.823e-18
c3668 n965__i1__i14__net1 vss 193.091e-18
c3669 n966__i1__i14__net1 vss 201.632e-18
c3670 n968__i1__i14__net1 vss 187.318e-18
c3671 n969__i1__i14__net1 vss 202.216e-18
c3672 n971__i1__i14__net1 vss 242.868e-18
c3673 n38__shift vss 47.0485e-18
c3674 n1264__vddio vss 268.738e-18
c3675 n1267__vddio vss 254.868e-18
c3676 n1268__vddio vss 134.679e-18
c3677 n1270__vddio vss 242.925e-18
c3678 n1271__vddio vss 139.901e-18
c3679 n1273__vddio vss 252.742e-18
c3680 n1274__vddio vss 137.738e-18
c3681 n1276__vddio vss 160.618e-18
c3682 n17__i5__i8__net2 vss 58.0624e-18
c3683 n8__i5__i6__net34 vss 130.538e-18
c3684 n912__i1__i14__net1 vss 229.933e-18
c3685 n914__i1__i14__net1 vss 196.891e-18
c3686 n915__i1__i14__net1 vss 236.092e-18
c3687 n917__i1__i14__net1 vss 274.512e-18
c3688 n920__i1__i14__net1 vss 229.252e-18
c3689 n923__i1__i14__net1 vss 194.615e-18
c3690 n924__i1__i14__net1 vss 219.939e-18
c3691 n926__i1__i14__net1 vss 196.852e-18
c3692 n927__i1__i14__net1 vss 206.757e-18
c3693 n929__i1__i14__net1 vss 190.044e-18
c3694 n930__i1__i14__net1 vss 205.891e-18
c3695 n932__i1__i14__net1 vss 244.793e-18
c3696 n27__i5__i8__net2 vss 193.113e-18
c3697 n109__i1__net2 vss 35.737e-18
c3698 n110__i1__net2 vss 47.715e-18
c3699 n35__shift vss 60.9169e-18
c3700 n1243__vddio vss 264.759e-18
c3701 n1244__vddio vss 252.682e-18
c3702 n1247__vddio vss 134.094e-18
c3703 n1248__vddio vss 240.386e-18
c3704 n1251__vddio vss 139.184e-18
c3705 n1252__vddio vss 251.592e-18
c3706 n1255__vddio vss 137.993e-18
c3707 n1262__vddio vss 162.119e-18
c3708 n54__reset vss 59.4144e-18
c3709 n97__i1__net2 vss 39.2353e-18
c3710 n98__i1__net2 vss 37.7237e-18
c3711 n2__i5__i6__net34 vss 117.838e-18
c3712 n872__i1__i14__net1 vss 135.109e-18
c3713 n873__i1__i14__net1 vss 213.779e-18
c3714 n875__i1__i14__net1 vss 196.891e-18
c3715 n876__i1__i14__net1 vss 219.887e-18
c3716 n878__i1__i14__net1 vss 256.004e-18
c3717 n881__i1__i14__net1 vss 256.508e-18
c3718 n884__i1__i14__net1 vss 182.256e-18
c3719 n885__i1__i14__net1 vss 207.184e-18
c3720 n887__i1__i14__net1 vss 184.192e-18
c3721 n888__i1__i14__net1 vss 226.811e-18
c3722 n890__i1__i14__net1 vss 178.134e-18
c3723 n891__i1__i14__net1 vss 227.193e-18
c3724 n893__i1__i14__net1 vss 233.763e-18
c3725 n7__i5__i8__i9__net24 vss 67.5198e-18
c3726 n6__i5__i8__i9__net23 vss 84.3725e-18
c3727 n89__i1__net2 vss 42.4364e-18
c3728 n90__i1__net2 vss 38.8751e-18
c3729 n198__vdd vss 88.2845e-18
c3730 n1222__vddio vss 286.649e-18
c3731 n1225__vddio vss 238.386e-18
c3732 n1226__vddio vss 151.358e-18
c3733 n1228__vddio vss 258.886e-18
c3734 n1229__vddio vss 156.638e-18
c3735 n1231__vddio vss 237.607e-18
c3736 n1232__vddio vss 155.355e-18
c3737 n1234__vddio vss 164.92e-18
c3738 n63__i5__clk_buf vss 114.8e-18
c3739 n6__i5__i8__i9__net24 vss 109.564e-18
c3740 n3__i5__i8__i9__net23 vss 97.9446e-18
c3741 n833__i1__i14__net1 vss 134.708e-18
c3742 n834__i1__i14__net1 vss 227.822e-18
c3743 n836__i1__i14__net1 vss 196.115e-18
c3744 n837__i1__i14__net1 vss 233.179e-18
c3745 n839__i1__i14__net1 vss 274.244e-18
c3746 n842__i1__i14__net1 vss 230.267e-18
c3747 n845__i1__i14__net1 vss 194.664e-18
c3748 n846__i1__i14__net1 vss 218.596e-18
c3749 n848__i1__i14__net1 vss 196.673e-18
c3750 n849__i1__i14__net1 vss 205.482e-18
c3751 n851__i1__i14__net1 vss 190.902e-18
c3752 n852__i1__i14__net1 vss 209.332e-18
c3753 n854__i1__i14__net1 vss 256.829e-18
c3754 n9__i5__i6__i4__net24 vss 57.8731e-18
c3755 n6__i5__i6__i4__net23 vss 82.5454e-18
c3756 n77__i1__net2 vss 29.0349e-18
c3757 n78__i1__net2 vss 38.3164e-18
c3758 n3__i5__i8__i9__net24 vss 106.815e-18
c3759 n2__i5__i8__i9__net23 vss 107.785e-18
c3760 n1201__vddio vss 271.48e-18
c3761 n1204__vddio vss 257.779e-18
c3762 n1205__vddio vss 136.358e-18
c3763 n1207__vddio vss 245.962e-18
c3764 n1208__vddio vss 141.61e-18
c3765 n1210__vddio vss 256.327e-18
c3766 n1211__vddio vss 140.274e-18
c3767 n1213__vddio vss 187.387e-18
c3768 n58__i5__clk_buf vss 119.821e-18
c3769 n6__i5__i6__i4__net24 vss 110.659e-18
c3770 n3__i5__i6__i4__net23 vss 98.2305e-18
c3771 n69__i1__net2 vss 39.1175e-18
c3772 n70__i1__net2 vss 46.7735e-18
c3773 n9__i5__i8__i9__net25 vss 110.709e-18
c3774 n6__i5__i8__i9__net21 vss 107.843e-18
c3775 n794__i1__i14__net1 vss 133.748e-18
c3776 n795__i1__i14__net1 vss 233.11e-18
c3777 n797__i1__i14__net1 vss 200.413e-18
c3778 n798__i1__i14__net1 vss 238.571e-18
c3779 n800__i1__i14__net1 vss 277.975e-18
c3780 n803__i1__i14__net1 vss 227.02e-18
c3781 n806__i1__i14__net1 vss 196.027e-18
c3782 n807__i1__i14__net1 vss 220.105e-18
c3783 n809__i1__i14__net1 vss 198.174e-18
c3784 n810__i1__i14__net1 vss 202.713e-18
c3785 n812__i1__i14__net1 vss 192.345e-18
c3786 n813__i1__i14__net1 vss 203.282e-18
c3787 n815__i1__i14__net1 vss 248.023e-18
c3788 n61__i1__net2 vss 30.8048e-18
c3789 n62__i1__net2 vss 58.4445e-18
c3790 n3__i5__i6__i4__net24 vss 107.133e-18
c3791 n2__i5__i6__i4__net23 vss 105.277e-18
c3792 n15__i5__i8__net4 vss 138.279e-18
c3793 n56__i5__clk_buf vss 152.88e-18
c3794 n6__i5__i8__i9__net25 vss 130.705e-18
c3795 n3__i5__i8__i9__net21 vss 88.8559e-18
c3796 n1174__vddio vss 142.291e-18
c3797 n1177__vddio vss 148.345e-18
c3798 n1178__vddio vss 72.0028e-18
c3799 n1180__vddio vss 131.286e-18
c3800 n1181__vddio vss 74.4314e-18
c3801 n1183__vddio vss 145.606e-18
c3802 n1184__vddio vss 73.0869e-18
c3803 n1186__vddio vss 143.772e-18
c3804 n9__i5__i8__net1 vss 50.1416e-18
c3805 n9__i5__i6__i4__net25 vss 101.765e-18
c3806 n6__i5__i6__i4__net21 vss 108.465e-18
c3807 n3__i5__i8__i9__net25 vss 90.5227e-18
c3808 n2__i5__i8__i9__net21 vss 112.785e-18
c3809 n29__i5__i6__net31 vss 116.403e-18
c3810 n51__i5__clk_buf vss 138.685e-18
c3811 n6__i5__i6__i4__net25 vss 114.351e-18
c3812 n3__i5__i6__i4__net21 vss 88.5725e-18
c3813 n12__i5__i8__net4 vss 130.421e-18
c3814 n3__i5__i6__i4__net25 vss 81.73e-18
c3815 n2__i5__i6__i4__net21 vss 94.4736e-18
c3816 n15__i5__i6__net33 vss 66.827e-18
c3817 n9__i5__i6__net33 vss 57.8082e-18
c3818 n44__i5__clk_buf vss 45.1627e-18
c3819 n11__i5__r1 vss 96.0145e-18
c3820 n159__vdd vss 54.3316e-18
c3821 n160__vdd vss 72.5992e-18
c3822 n28__shift vss 44.1594e-18
c3823 n158__vdd vss 8.51146e-18
c3824 n8__i5__i6__net32 vss 129.536e-18
c3825 n1100__vddio vss 146.312e-18
c3826 n1103__vddio vss 134.718e-18
c3827 n1104__vddio vss 73.9053e-18
c3828 n1106__vddio vss 132.666e-18
c3829 n1107__vddio vss 76.7107e-18
c3830 n1109__vddio vss 136.733e-18
c3831 n1110__vddio vss 76.5474e-18
c3832 n1112__vddio vss 117.273e-18
c3833 n157__vdd vss 57.2499e-18
c3834 n773__i1__i14__net1 vss 51.3611e-18
c3835 n774__i1__i14__net1 vss 44.7569e-18
c3836 n1909__chipdriverout vss 222.882e-18
c3837 n1911__chipdriverout vss 192.29e-18
c3838 n1912__chipdriverout vss 228.128e-18
c3839 n1914__chipdriverout vss 269.027e-18
c3840 n1891__chipdriverout vss 232.68e-18
c3841 n1894__chipdriverout vss 203.171e-18
c3842 n1895__chipdriverout vss 229.258e-18
c3843 n1897__chipdriverout vss 205.374e-18
c3844 n1898__chipdriverout vss 211.39e-18
c3845 n1900__chipdriverout vss 199.048e-18
c3846 n1901__chipdriverout vss 211.691e-18
c3847 n1903__chipdriverout vss 255.192e-18
c3848 n154__vdd vss 63.7987e-18
c3849 n151__vdd vss 46.2891e-18
c3850 n22__shift vss 61.2388e-18
c3851 n769__i1__i14__net1 vss 36.2924e-18
c3852 n770__i1__i14__net1 vss 46.0224e-18
c3853 n1079__vddio vss 264.419e-18
c3854 n1082__vddio vss 252.613e-18
c3855 n1083__vddio vss 134.138e-18
c3856 n1085__vddio vss 240.454e-18
c3857 n1086__vddio vss 139.162e-18
c3858 n1088__vddio vss 251.765e-18
c3859 n1089__vddio vss 138.102e-18
c3860 n1091__vddio vss 162.355e-18
c3861 n765__i1__i14__net1 vss 39.1199e-18
c3862 n766__i1__i14__net1 vss 47.6055e-18
c3863 n2__i5__i6__net32 vss 117.595e-18
c3864 n1869__chipdriverout vss 130.998e-18
c3865 n1870__chipdriverout vss 220.999e-18
c3866 n1872__chipdriverout vss 190.226e-18
c3867 n1873__chipdriverout vss 226.466e-18
c3868 n1875__chipdriverout vss 264.048e-18
c3869 n1852__chipdriverout vss 237.422e-18
c3870 n1855__chipdriverout vss 203.697e-18
c3871 n1856__chipdriverout vss 230.761e-18
c3872 n1858__chipdriverout vss 206.051e-18
c3873 n1859__chipdriverout vss 217.635e-18
c3874 n1861__chipdriverout vss 199.602e-18
c3875 n1862__chipdriverout vss 218.253e-18
c3876 n1864__chipdriverout vss 258.693e-18
c3877 n8__clk_out vss 68.7481e-18
c3878 n1058__vddio vss 282.096e-18
c3879 n1061__vddio vss 248.859e-18
c3880 n1062__vddio vss 156.133e-18
c3881 n1064__vddio vss 269.263e-18
c3882 n1065__vddio vss 161.826e-18
c3883 n1067__vddio vss 247.325e-18
c3884 n1068__vddio vss 160.12e-18
c3885 n1070__vddio vss 196.687e-18
c3886 n40__reset vss 62.0992e-18
c3887 n9__i5__r2 vss 71.4816e-18
c3888 n1829__chipdriverout vss 258.524e-18
c3889 n1832__chipdriverout vss 197.34e-18
c3890 n1833__chipdriverout vss 222.427e-18
c3891 n1835__chipdriverout vss 199.315e-18
c3892 n1836__chipdriverout vss 225.717e-18
c3893 n1838__chipdriverout vss 177.437e-18
c3894 n1839__chipdriverout vss 225.808e-18
c3895 n1841__chipdriverout vss 252.185e-18
c3896 n1812__chipdriverout vss 126.312e-18
c3897 n1815__chipdriverout vss 200.558e-18
c3898 n1816__chipdriverout vss 185.752e-18
c3899 n1819__chipdriverout vss 221.343e-18
c3900 n1820__chipdriverout vss 264.103e-18
c3901 n9__i5__i6__i2__net24 vss 57.9076e-18
c3902 n6__i5__i6__i2__net23 vss 81.0036e-18
c3903 n753__i1__i14__net1 vss 43.627e-18
c3904 n754__i1__i14__net1 vss 36.4915e-18
c3905 n1037__vddio vss 270.982e-18
c3906 n1040__vddio vss 238.063e-18
c3907 n1041__vddio vss 150.913e-18
c3908 n1043__vddio vss 258.962e-18
c3909 n1044__vddio vss 156.136e-18
c3910 n1046__vddio vss 236.375e-18
c3911 n1047__vddio vss 154.838e-18
c3912 n1049__vddio vss 162.545e-18
c3913 n35__i5__clk_buf vss 120.604e-18
c3914 n6__i5__i6__i2__net24 vss 110.503e-18
c3915 n3__i5__i6__i2__net23 vss 98.983e-18
c3916 n749__i1__i14__net1 vss 39.2398e-18
c3917 n750__i1__i14__net1 vss 34.2851e-18
c3918 n1791__chipdriverout vss 144.043e-18
c3919 n1792__chipdriverout vss 201.996e-18
c3920 n1794__chipdriverout vss 170.962e-18
c3921 n1795__chipdriverout vss 206.791e-18
c3922 n1797__chipdriverout vss 245.009e-18
c3923 n1774__chipdriverout vss 254.08e-18
c3924 n1777__chipdriverout vss 180.1e-18
c3925 n1778__chipdriverout vss 205.149e-18
c3926 n1780__chipdriverout vss 182.002e-18
c3927 n1781__chipdriverout vss 224.506e-18
c3928 n1783__chipdriverout vss 176.032e-18
c3929 n1784__chipdriverout vss 224.59e-18
c3930 n1786__chipdriverout vss 230.374e-18
c3931 n8__i5__i7__i7__net3 vss 119.006e-18
c3932 n3__i5__i6__i2__net24 vss 107.849e-18
c3933 n2__i5__i6__i2__net23 vss 105.919e-18
c3934 n745__i1__i14__net1 vss 35.7003e-18
c3935 n746__i1__i14__net1 vss 44.1487e-18
c3936 n1005__vddio vss 278.416e-18
c3937 n1008__vddio vss 229.86e-18
c3938 n1009__vddio vss 146.532e-18
c3939 n1012__vddio vss 250.187e-18
c3940 n1013__vddio vss 151.585e-18
c3941 n1016__vddio vss 228.843e-18
c3942 n1017__vddio vss 149.403e-18
c3943 n1025__vddio vss 178.273e-18
c3944 n27__i5__i7__i7__net1 vss 145.32e-18
c3945 n9__i5__i6__i2__net25 vss 101.357e-18
c3946 n6__i5__i6__i2__net21 vss 107.323e-18
c3947 n741__i1__i14__net1 vss 46.4724e-18
c3948 n742__i1__i14__net1 vss 47.4103e-18
c3949 n23__i5__i7__net46 vss 156.545e-18
c3950 n1752__chipdriverout vss 127.911e-18
c3951 n1753__chipdriverout vss 218.187e-18
c3952 n1755__chipdriverout vss 187.412e-18
c3953 n1756__chipdriverout vss 223.329e-18
c3954 n1758__chipdriverout vss 264.158e-18
c3955 n1735__chipdriverout vss 233.986e-18
c3956 n1738__chipdriverout vss 199.118e-18
c3957 n1739__chipdriverout vss 224.992e-18
c3958 n1741__chipdriverout vss 201.235e-18
c3959 n1742__chipdriverout vss 212.094e-18
c3960 n1744__chipdriverout vss 194.707e-18
c3961 n1745__chipdriverout vss 211.396e-18
c3962 n1747__chipdriverout vss 249.719e-18
c3963 n17__i5__i6__net31 vss 117.107e-18
c3964 n1555__vddio vss 6.62809e-18
c3965 n737__i1__i14__net1 vss 43.7208e-18
c3966 n738__i1__i14__net1 vss 37.2656e-18
c3967 n6__i5__i6__i2__net25 vss 113.987e-18
c3968 n3__i5__i6__i2__net21 vss 87.978e-18
c3969 n985__vddio vss 281.515e-18
c3970 n988__vddio vss 235.237e-18
c3971 n989__vddio vss 149.528e-18
c3972 n991__vddio vss 255.576e-18
c3973 n992__vddio vss 154.698e-18
c3974 n994__vddio vss 234.117e-18
c3975 n995__vddio vss 153.369e-18
c3976 n997__vddio vss 185.404e-18
c3977 n18__i5__i7__net46 vss 138.334e-18
c3978 n733__i1__i14__net1 vss 46.49e-18
c3979 n734__i1__i14__net1 vss 38.6591e-18
c3980 n3__i5__i6__i2__net25 vss 82.6089e-18
c3981 n2__i5__i6__i2__net21 vss 94.828e-18
c3982 n15__i5__i6__net30 vss 68.2143e-18
c3983 n1713__chipdriverout vss 16.7041e-18
c3984 n1714__chipdriverout vss 203.816e-18
c3985 n1716__chipdriverout vss 172.447e-18
c3986 n1717__chipdriverout vss 208.869e-18
c3987 n1719__chipdriverout vss 245.586e-18
c3988 n1696__chipdriverout vss 259.764e-18
c3989 n1699__chipdriverout vss 186.625e-18
c3990 n1700__chipdriverout vss 212.619e-18
c3991 n1702__chipdriverout vss 188.622e-18
c3992 n1703__chipdriverout vss 232.06e-18
c3993 n1705__chipdriverout vss 182.53e-18
c3994 n1706__chipdriverout vss 232.601e-18
c3995 n1708__chipdriverout vss 239.763e-18
c3996 n729__i1__i14__net1 vss 43.7208e-18
c3997 n730__i1__i14__net1 vss 38.4099e-18
c3998 n21__i5__i7__net44 vss 122.478e-18
c3999 n9__i5__i6__net30 vss 58.3495e-18
c4000 n964__vddio vss 274.882e-18
c4001 n967__vddio vss 262.932e-18
c4002 n968__vddio vss 139.482e-18
c4003 n970__vddio vss 251.093e-18
c4004 n971__vddio vss 144.784e-18
c4005 n973__vddio vss 261.398e-18
c4006 n974__vddio vss 143.524e-18
c4007 n976__vddio vss 167.984e-18
c4008 n4__i5__r2 vss 96.234e-18
c4009 n725__i1__i14__net1 vss 39.2159e-18
c4010 n726__i1__i14__net1 vss 47.5829e-18
c4011 n1675__chipdriverout vss 218.23e-18
c4012 n1677__chipdriverout vss 188.069e-18
c4013 n1678__chipdriverout vss 223.408e-18
c4014 n1680__chipdriverout vss 263.189e-18
c4015 n1657__chipdriverout vss 233.641e-18
c4016 n1660__chipdriverout vss 198.664e-18
c4017 n1661__chipdriverout vss 224.661e-18
c4018 n1663__chipdriverout vss 200.862e-18
c4019 n1664__chipdriverout vss 211.696e-18
c4020 n1666__chipdriverout vss 194.55e-18
c4021 n1667__chipdriverout vss 211.989e-18
c4022 n1669__chipdriverout vss 248.773e-18
c4023 n721__i1__i14__net1 vss 35.7412e-18
c4024 n722__i1__i14__net1 vss 45.5269e-18
c4025 n47__vdd vss 109.101e-18
c4026 n15__shift vss 38.731e-18
c4027 n943__vddio vss 287.252e-18
c4028 n946__vddio vss 240.748e-18
c4029 n947__vddio vss 152.077e-18
c4030 n949__vddio vss 261.403e-18
c4031 n950__vddio vss 157.453e-18
c4032 n952__vddio vss 239.06e-18
c4033 n953__vddio vss 156.003e-18
c4034 n955__vddio vss 163.845e-18
c4035 n44__vdd vss 99.6706e-18
c4036 n717__i1__i14__net1 vss 46.7265e-18
c4037 n718__i1__i14__net1 vss 38.5804e-18
c4038 n46__vdd vss 63.9379e-18
c4039 n1635__chipdriverout vss 133.375e-18
c4040 n1636__chipdriverout vss 223.722e-18
c4041 n1638__chipdriverout vss 191.957e-18
c4042 n1639__chipdriverout vss 229.113e-18
c4043 n1641__chipdriverout vss 266.915e-18
c4044 n1618__chipdriverout vss 234.344e-18
c4045 n1621__chipdriverout vss 199.751e-18
c4046 n1622__chipdriverout vss 226.191e-18
c4047 n1624__chipdriverout vss 202.035e-18
c4048 n1625__chipdriverout vss 213.114e-18
c4049 n1627__chipdriverout vss 195.501e-18
c4050 n1628__chipdriverout vss 213.522e-18
c4051 n1630__chipdriverout vss 253.714e-18
c4052 n21__i5__i7__i7__net1 vss 79.929e-18
c4053 n709__i1__i14__net1 vss 37.3472e-18
c4054 n710__i1__i14__net1 vss 45.5112e-18
c4055 n9__shift vss 62.0944e-18
c4056 n922__vddio vss 267.687e-18
c4057 n925__vddio vss 252.994e-18
c4058 n926__vddio vss 133.234e-18
c4059 n928__vddio vss 240.876e-18
c4060 n929__vddio vss 139.266e-18
c4061 n931__vddio vss 252.618e-18
c4062 n932__vddio vss 137.657e-18
c4063 n934__vddio vss 160.331e-18
c4064 n12__i5__i6__net31 vss 15.5277e-18
c4065 n1581__chipdriverout vss 135.109e-18
c4066 n1582__chipdriverout vss 229.932e-18
c4067 n1584__chipdriverout vss 196.861e-18
c4068 n1585__chipdriverout vss 235.352e-18
c4069 n1587__chipdriverout vss 273.178e-18
c4070 n1590__chipdriverout vss 236.098e-18
c4071 n1593__chipdriverout vss 200.663e-18
c4072 n1594__chipdriverout vss 225.602e-18
c4073 n1596__chipdriverout vss 202.651e-18
c4074 n1597__chipdriverout vss 213.539e-18
c4075 n1599__chipdriverout vss 197.308e-18
c4076 n1600__chipdriverout vss 214.133e-18
c4077 n1602__chipdriverout vss 252.373e-18
c4078 n1559__vddio vss 7.25738e-18
c4079 n693__i1__i14__net1 vss 42.611e-18
c4080 n694__i1__i14__net1 vss 38.5043e-18
c4081 n891__vddio vss 270.873e-18
c4082 n894__vddio vss 238.163e-18
c4083 n895__vddio vss 150.371e-18
c4084 n897__vddio vss 258.531e-18
c4085 n898__vddio vss 156.394e-18
c4086 n900__vddio vss 237.728e-18
c4087 n901__vddio vss 154.359e-18
c4088 n903__vddio vss 184.794e-18
c4089 n3__i5__r1 vss 85.1055e-18
c4090 n5__i5__r1 vss 56.027e-18
c4091 n1541__chipdriverout vss 135.958e-18
c4092 n1542__chipdriverout vss 231.367e-18
c4093 n1544__chipdriverout vss 197.279e-18
c4094 n1545__chipdriverout vss 237.121e-18
c4095 n1547__chipdriverout vss 273.238e-18
c4096 n1550__chipdriverout vss 231.336e-18
c4097 n1553__chipdriverout vss 196.43e-18
c4098 n1554__chipdriverout vss 221.361e-18
c4099 n1556__chipdriverout vss 198.506e-18
c4100 n1557__chipdriverout vss 209.227e-18
c4101 n1559__chipdriverout vss 192.94e-18
c4102 n1560__chipdriverout vss 209.252e-18
c4103 n1562__chipdriverout vss 247.772e-18
c4104 n17__i5__clk_buf vss 41.6988e-18
c4105 n13__i5__i7__net46 vss 117.647e-18
c4106 n19__i5__i7__i7__net1 vss 240.844e-18
c4107 n870__vddio vss 251.864e-18
c4108 n871__vddio vss 252.437e-18
c4109 n874__vddio vss 133.312e-18
c4110 n875__vddio vss 240.483e-18
c4111 n878__vddio vss 139.194e-18
c4112 n879__vddio vss 251.389e-18
c4113 n882__vddio vss 136.864e-18
c4114 n889__vddio vss 159.619e-18
c4115 n12__i5__i7__i6__net1 vss 117.313e-18
c4116 n1501__chipdriverout vss 151.349e-18
c4117 n1502__chipdriverout vss 229.962e-18
c4118 n1504__chipdriverout vss 180.479e-18
c4119 n1505__chipdriverout vss 235.382e-18
c4120 n1507__chipdriverout vss 273.209e-18
c4121 n1510__chipdriverout vss 221.04e-18
c4122 n1513__chipdriverout vss 186.632e-18
c4123 n1514__chipdriverout vss 209.882e-18
c4124 n1516__chipdriverout vss 188.773e-18
c4125 n1517__chipdriverout vss 197.01e-18
c4126 n1519__chipdriverout vss 183.098e-18
c4127 n1520__chipdriverout vss 197.75e-18
c4128 n1522__chipdriverout vss 238.273e-18
c4129 n6__i5__r0 vss 98.5681e-18
c4130 n8__i5__r0 vss 95.2444e-18
c4131 n661__i1__i14__net1 vss 42.611e-18
c4132 n662__i1__i14__net1 vss 38.6706e-18
c4133 n16__i5__i7__i7__net1 vss 91.9313e-18
c4134 n849__vddio vss 270.162e-18
c4135 n852__vddio vss 255.8e-18
c4136 n853__vddio vss 135.381e-18
c4137 n855__vddio vss 243.979e-18
c4138 n856__vddio vss 141.151e-18
c4139 n858__vddio vss 255.468e-18
c4140 n859__vddio vss 139.854e-18
c4141 n861__vddio vss 186.916e-18
c4142 n653__i1__i14__net1 vss 46.8202e-18
c4143 n654__i1__i14__net1 vss 37.5286e-18
c4144 n1447__chipdriverout vss 229.194e-18
c4145 n1450__chipdriverout vss 180.158e-18
c4146 n1451__chipdriverout vss 234.564e-18
c4147 n1454__chipdriverout vss 253.971e-18
c4148 n1455__chipdriverout vss 246.207e-18
c4149 n1458__chipdriverout vss 174.57e-18
c4150 n1459__chipdriverout vss 213.263e-18
c4151 n1462__chipdriverout vss 176.456e-18
c4152 n1463__chipdriverout vss 216.449e-18
c4153 n1466__chipdriverout vss 171.047e-18
c4154 n1467__chipdriverout vss 217.358e-18
c4155 n1470__chipdriverout vss 226.296e-18
c4156 n17__i5__i7__net50 vss 166.622e-18
c4157 n828__vddio vss 273.197e-18
c4158 n829__vddio vss 256.245e-18
c4159 n832__vddio vss 136.654e-18
c4160 n833__vddio vss 245.954e-18
c4161 n836__vddio vss 141.85e-18
c4162 n837__vddio vss 256.245e-18
c4163 n840__vddio vss 140.63e-18
c4164 n847__vddio vss 166.178e-18
c4165 n15__i5__i7__net50 vss 145.615e-18
c4166 n18__i5__i7__net51 vss 104.582e-18
c4167 n633__i1__i14__net1 vss 45.7602e-18
c4168 n634__i1__i14__net1 vss 38.3303e-18
c4169 n12__i5__i7__net44 vss 71.5025e-18
c4170 n1407__chipdriverout vss 150.112e-18
c4171 n1408__chipdriverout vss 212.548e-18
c4172 n1410__chipdriverout vss 179.999e-18
c4173 n1411__chipdriverout vss 217.682e-18
c4174 n1413__chipdriverout vss 253.018e-18
c4175 n1416__chipdriverout vss 256.083e-18
c4176 n1419__chipdriverout vss 184.379e-18
c4177 n1420__chipdriverout vss 208.898e-18
c4178 n1422__chipdriverout vss 186.204e-18
c4179 n1423__chipdriverout vss 227.864e-18
c4180 n1425__chipdriverout vss 180.682e-18
c4181 n1426__chipdriverout vss 233.125e-18
c4182 n1428__chipdriverout vss 234.611e-18
c4183 n4__i5__i7__net46 vss 147.143e-18
c4184 n625__i1__i14__net1 vss 42.7048e-18
c4185 n626__i1__i14__net1 vss 38.5406e-18
c4186 n11__i5__i7__i7__net1 vss 66.5637e-18
c4187 n13__i5__i7__i7__net1 vss 47.3398e-18
c4188 n801__vddio vss 285.159e-18
c4189 n804__vddio vss 238.163e-18
c4190 n805__vddio vss 150.371e-18
c4191 n807__vddio vss 258.531e-18
c4192 n808__vddio vss 156.394e-18
c4193 n810__vddio vss 237.833e-18
c4194 n811__vddio vss 154.848e-18
c4195 n813__vddio vss 185.644e-18
c4196 n9__i5__i7__net50 vss 145.214e-18
c4197 n621__i1__i14__net1 vss 46.7264e-18
c4198 n622__i1__i14__net1 vss 36.8186e-18
c4199 n9__i5__i7__net44 vss 174.334e-18
c4200 n1368__chipdriverout vss 151.803e-18
c4201 n1369__chipdriverout vss 213.866e-18
c4202 n1371__chipdriverout vss 196.775e-18
c4203 n1372__chipdriverout vss 219.066e-18
c4204 n1374__chipdriverout vss 273.239e-18
c4205 n1377__chipdriverout vss 231.3e-18
c4206 n1380__chipdriverout vss 196.331e-18
c4207 n1381__chipdriverout vss 204.997e-18
c4208 n1383__chipdriverout vss 198.392e-18
c4209 n1384__chipdriverout vss 209.104e-18
c4210 n1386__chipdriverout vss 193.116e-18
c4211 n1387__chipdriverout vss 209.89e-18
c4212 n1389__chipdriverout vss 248.499e-18
c4213 n12__i5__i7__net47 vss 165.505e-18
c4214 n613__i1__i14__net1 vss 35.7413e-18
c4215 n614__i1__i14__net1 vss 38.5406e-18
c4216 n776__vddio vss 279.611e-18
c4217 n779__vddio vss 231.704e-18
c4218 n780__vddio vss 146.122e-18
c4219 n782__vddio vss 251.714e-18
c4220 n783__vddio vss 152.26e-18
c4221 n785__vddio vss 231.245e-18
c4222 n786__vddio vss 150.328e-18
c4223 n788__vddio vss 178.624e-18
c4224 n601__i1__i14__net1 vss 38.1504e-18
c4225 n602__i1__i14__net1 vss 42.3214e-18
c4226 n1329__chipdriverout vss 129.023e-18
c4227 n1330__chipdriverout vss 203.379e-18
c4228 n1332__chipdriverout vss 188.467e-18
c4229 n1333__chipdriverout vss 208.042e-18
c4230 n1335__chipdriverout vss 249.309e-18
c4231 n1338__chipdriverout vss 248.619e-18
c4232 n1341__chipdriverout vss 173.623e-18
c4233 n1342__chipdriverout vss 196.713e-18
c4234 n1344__chipdriverout vss 175.471e-18
c4235 n1345__chipdriverout vss 216.753e-18
c4236 n1347__chipdriverout vss 170.559e-18
c4237 n1348__chipdriverout vss 216.446e-18
c4238 n1350__chipdriverout vss 223.341e-18
c4239 n10__i5__i7__net47 vss 97.3053e-18
c4240 n15__i5__i7__net51 vss 98.4801e-18
c4241 n597__i1__i14__net1 vss 45.7283e-18
c4242 n598__i1__i14__net1 vss 26.1498e-18
c4243 n755__vddio vss 270.367e-18
c4244 n758__vddio vss 235.89e-18
c4245 n759__vddio vss 149.28e-18
c4246 n761__vddio vss 256.425e-18
c4247 n762__vddio vss 155.284e-18
c4248 n764__vddio vss 235.342e-18
c4249 n765__vddio vss 152.4e-18
c4250 n767__vddio vss 160.225e-18
c4251 n1290__chipdriverout vss 129.346e-18
c4252 n1291__chipdriverout vss 219.774e-18
c4253 n1293__chipdriverout vss 188.848e-18
c4254 n1294__chipdriverout vss 225.043e-18
c4255 n1296__chipdriverout vss 264.166e-18
c4256 n1299__chipdriverout vss 234.323e-18
c4257 n1302__chipdriverout vss 200.044e-18
c4258 n1303__chipdriverout vss 226.065e-18
c4259 n1305__chipdriverout vss 202.416e-18
c4260 n1306__chipdriverout vss 213.356e-18
c4261 n1308__chipdriverout vss 196.708e-18
c4262 n1309__chipdriverout vss 214.041e-18
c4263 n1311__chipdriverout vss 253.914e-18
c4264 n581__i1__i14__net1 vss 46.6387e-18
c4265 n582__i1__i14__net1 vss 26.03e-18
c4266 n734__vddio vss 279.82e-18
c4267 n737__vddio vss 247.251e-18
c4268 n738__vddio vss 155.674e-18
c4269 n740__vddio vss 267.88e-18
c4270 n741__vddio vss 161.648e-18
c4271 n743__vddio vss 246.478e-18
c4272 n744__vddio vss 160.052e-18
c4273 n746__vddio vss 191.385e-18
c4274 n12__i5__i7__i5__net1 vss 117.605e-18
c4275 n12__i5__i7__i4__net1 vss 117.807e-18
c4276 n573__i1__i14__net1 vss 36.4245e-18
c4277 n574__i1__i14__net1 vss 47.6925e-18
c4278 n10__i5__i7__net51 vss 126.979e-18
c4279 n12__i5__i7__net51 vss 97.8632e-18
c4280 n6__i5__i7__net50 vss 153.704e-18
c4281 n8__i5__i7__net50 vss 95.0585e-18
c4282 n1251__chipdriverout vss 145.737e-18
c4283 n1252__chipdriverout vss 219.184e-18
c4284 n1254__chipdriverout vss 188.254e-18
c4285 n1255__chipdriverout vss 208.525e-18
c4286 n1257__chipdriverout vss 243.111e-18
c4287 n1260__chipdriverout vss 261.799e-18
c4288 n1263__chipdriverout vss 188.198e-18
c4289 n1264__chipdriverout vss 214.232e-18
c4290 n1266__chipdriverout vss 190.216e-18
c4291 n1267__chipdriverout vss 233.782e-18
c4292 n1269__chipdriverout vss 184.101e-18
c4293 n1270__chipdriverout vss 234.337e-18
c4294 n1272__chipdriverout vss 241.253e-18
c4295 n565__i1__i14__net1 vss 38.5181e-18
c4296 n566__i1__i14__net1 vss 47.4842e-18
c4297 n713__vddio vss 267.492e-18
c4298 n716__vddio vss 255.958e-18
c4299 n717__vddio vss 135.676e-18
c4300 n719__vddio vss 243.566e-18
c4301 n720__vddio vss 140.892e-18
c4302 n722__vddio vss 255.111e-18
c4303 n723__vddio vss 139.637e-18
c4304 n725__vddio vss 163.879e-18
c4305 n17__i5__i7__xor3 vss 168.214e-18
c4306 n17__i5__i7__xor0 vss 164.369e-18
c4307 n557__i1__i14__net1 vss 36.5298e-18
c4308 n558__i1__i14__net1 vss 46.9698e-18
c4309 n1213__chipdriverout vss 217.638e-18
c4310 n1215__chipdriverout vss 187.337e-18
c4311 n1216__chipdriverout vss 222.849e-18
c4312 n1218__chipdriverout vss 262.572e-18
c4313 n1221__chipdriverout vss 233.149e-18
c4314 n1224__chipdriverout vss 198.14e-18
c4315 n1225__chipdriverout vss 223.476e-18
c4316 n1227__chipdriverout vss 200.278e-18
c4317 n1228__chipdriverout vss 210.405e-18
c4318 n1230__chipdriverout vss 194.018e-18
c4319 n1231__chipdriverout vss 210.566e-18
c4320 n1233__chipdriverout vss 256.022e-18
c4321 n15__i5__i7__xor3 vss 148.42e-18
c4322 n15__i5__i7__xor0 vss 100.048e-18
c4323 n549__i1__i14__net1 vss 45.6596e-18
c4324 n550__i1__i14__net1 vss 47.4216e-18
c4325 n18__i5__i7__xor2 vss 83.6383e-18
c4326 n19__i5__i7__xor1 vss 103.024e-18
c4327 n692__vddio vss 263.304e-18
c4328 n695__vddio vss 249.592e-18
c4329 n696__vddio vss 132.101e-18
c4330 n698__vddio vss 237.066e-18
c4331 n699__vddio vss 137.196e-18
c4332 n701__vddio vss 248.73e-18
c4333 n702__vddio vss 135.973e-18
c4334 n704__vddio vss 182.504e-18
c4335 n537__i1__i14__net1 vss 43.9192e-18
c4336 n538__i1__i14__net1 vss 36.2633e-18
c4337 n7__i5__i7__net47 vss 150.265e-18
c4338 n4__i5__i7__net44 vss 81.4412e-18
c4339 n1173__chipdriverout vss 125.159e-18
c4340 n1174__chipdriverout vss 199.551e-18
c4341 n1176__chipdriverout vss 184.879e-18
c4342 n1177__chipdriverout vss 204.03e-18
c4343 n1179__chipdriverout vss 244.368e-18
c4344 n1182__chipdriverout vss 257.934e-18
c4345 n1185__chipdriverout vss 181.697e-18
c4346 n1186__chipdriverout vss 205.406e-18
c4347 n1188__chipdriverout vss 183.399e-18
c4348 n1189__chipdriverout vss 225.247e-18
c4349 n1191__chipdriverout vss 177.523e-18
c4350 n1192__chipdriverout vss 225.096e-18
c4351 n1194__chipdriverout vss 230.025e-18
c4352 n533__i1__i14__net1 vss 45.3323e-18
c4353 n534__i1__i14__net1 vss 27.8637e-18
c4354 n10__i5__i7__i5__net1 vss 226.176e-18
c4355 n10__i5__i7__i4__net1 vss 129.256e-18
c4356 n9__i5__i7__xor3 vss 148.855e-18
c4357 n9__i5__i7__xor0 vss 146.93e-18
c4358 n671__vddio vss 256.279e-18
c4359 n672__vddio vss 253.494e-18
c4360 n675__vddio vss 134.081e-18
c4361 n676__vddio vss 241.724e-18
c4362 n679__vddio vss 139.236e-18
c4363 n680__vddio vss 251.816e-18
c4364 n683__vddio vss 137.961e-18
c4365 n690__vddio vss 184.16e-18
c4366 n1134__chipdriverout vss 144.137e-18
c4367 n1135__chipdriverout vss 202.341e-18
c4368 n1137__chipdriverout vss 171.129e-18
c4369 n1138__chipdriverout vss 207.278e-18
c4370 n1140__chipdriverout vss 245.603e-18
c4371 n1143__chipdriverout vss 257.704e-18
c4372 n1146__chipdriverout vss 183.152e-18
c4373 n1147__chipdriverout vss 208.35e-18
c4374 n1149__chipdriverout vss 185.054e-18
c4375 n1150__chipdriverout vss 227.932e-18
c4376 n1152__chipdriverout vss 179.028e-18
c4377 n1153__chipdriverout vss 228.229e-18
c4378 n1155__chipdriverout vss 232.225e-18
c4379 n517__i1__i14__net1 vss 38.7599e-18
c4380 n518__i1__i14__net1 vss 36.0082e-18
c4381 n650__vddio vss 261.733e-18
c4382 n653__vddio vss 259.501e-18
c4383 n654__vddio vss 137.696e-18
c4384 n656__vddio vss 247.929e-18
c4385 n657__vddio vss 142.872e-18
c4386 n659__vddio vss 257.76e-18
c4387 n660__vddio vss 141.19e-18
c4388 n662__vddio vss 188.245e-18
c4389 n509__i1__i14__net1 vss 43.4248e-18
c4390 n510__i1__i14__net1 vss 38.2541e-18
c4391 n15__i5__i7__xor2 vss 125.371e-18
c4392 n15__i5__i7__xor1 vss 68.6008e-18
c4393 n1093__chipdriverout vss 147.91e-18
c4394 n1094__chipdriverout vss 206.187e-18
c4395 n1097__chipdriverout vss 174.304e-18
c4396 n1098__chipdriverout vss 211.534e-18
c4397 n1101__chipdriverout vss 245.653e-18
c4398 n1102__chipdriverout vss 260.231e-18
c4399 n1105__chipdriverout vss 187.86e-18
c4400 n1106__chipdriverout vss 214.485e-18
c4401 n1109__chipdriverout vss 190.006e-18
c4402 n1110__chipdriverout vss 233.721e-18
c4403 n1113__chipdriverout vss 183.666e-18
c4404 n1114__chipdriverout vss 233.261e-18
c4405 n1117__chipdriverout vss 241.876e-18
c4406 n501__i1__i14__net1 vss 38.7086e-18
c4407 n502__i1__i14__net1 vss 34.2752e-18
c4408 n619__vddio vss 256.517e-18
c4409 n622__vddio vss 258.407e-18
c4410 n623__vddio vss 136.837e-18
c4411 n625__vddio vss 245.906e-18
c4412 n626__vddio vss 142.192e-18
c4413 n628__vddio vss 256.952e-18
c4414 n629__vddio vss 140.323e-18
c4415 n631__vddio vss 163.979e-18
c4416 n489__i1__i14__net1 vss 43.8685e-18
c4417 n490__i1__i14__net1 vss 37.6103e-18
c4418 n1056__chipdriverout vss 147.46e-18
c4419 n1057__chipdriverout vss 202.828e-18
c4420 n1059__chipdriverout vss 171.612e-18
c4421 n1060__chipdriverout vss 207.772e-18
c4422 n1062__chipdriverout vss 244.375e-18
c4423 n1065__chipdriverout vss 256.241e-18
c4424 n1068__chipdriverout vss 182.146e-18
c4425 n1069__chipdriverout vss 207.037e-18
c4426 n1071__chipdriverout vss 184.067e-18
c4427 n1072__chipdriverout vss 226.621e-18
c4428 n1074__chipdriverout vss 178.082e-18
c4429 n1075__chipdriverout vss 227.14e-18
c4430 n1077__chipdriverout vss 234.767e-18
c4431 n485__i1__i14__net1 vss 38.1434e-18
c4432 n486__i1__i14__net1 vss 34.1087e-18
c4433 n598__vddio vss 250.841e-18
c4434 n599__vddio vss 252.507e-18
c4435 n602__vddio vss 133.984e-18
c4436 n603__vddio vss 240.164e-18
c4437 n606__vddio vss 139.058e-18
c4438 n607__vddio vss 251.686e-18
c4439 n610__vddio vss 137.945e-18
c4440 n617__vddio vss 162.147e-18
c4441 n6__i5__i7__xor3 vss 73.0273e-18
c4442 n8__i5__i7__xor3 vss 142.283e-18
c4443 n6__i5__i7__xor0 vss 72.8113e-18
c4444 n8__i5__i7__xor0 vss 147.829e-18
c4445 n473__i1__i14__net1 vss 44.9317e-18
c4446 n474__i1__i14__net1 vss 37.6103e-18
c4447 n1017__chipdriverout vss 128.862e-18
c4448 n1018__chipdriverout vss 210.89e-18
c4449 n1020__chipdriverout vss 194.565e-18
c4450 n1021__chipdriverout vss 215.876e-18
c4451 n1023__chipdriverout vss 256.937e-18
c4452 n1026__chipdriverout vss 252.91e-18
c4453 n1029__chipdriverout vss 177.27e-18
c4454 n1030__chipdriverout vss 200.64e-18
c4455 n1032__chipdriverout vss 178.884e-18
c4456 n1033__chipdriverout vss 220.56e-18
c4457 n1035__chipdriverout vss 173.13e-18
c4458 n1036__chipdriverout vss 220.312e-18
c4459 n1038__chipdriverout vss 224.94e-18
c4460 n13__i5__i7__x3out vss 112.397e-18
c4461 n13__i5__i7__x0out vss 121.809e-18
c4462 n14__i5__i7__y3out vss 139.31e-18
c4463 n16__i5__i7__y0out vss 186.989e-18
c4464 n577__vddio vss 255.754e-18
c4465 n580__vddio vss 253.293e-18
c4466 n581__vddio vss 134.548e-18
c4467 n583__vddio vss 241.793e-18
c4468 n584__vddio vss 139.485e-18
c4469 n586__vddio vss 251.932e-18
c4470 n587__vddio vss 138.524e-18
c4471 n589__vddio vss 163.467e-18
c4472 n461__i1__i14__net1 vss 42.1817e-18
c4473 n462__i1__i14__net1 vss 39.6514e-18
c4474 n976__chipdriverout vss 18.7842e-18
c4475 n977__chipdriverout vss 214.726e-18
c4476 n980__chipdriverout vss 181.546e-18
c4477 n981__chipdriverout vss 220.046e-18
c4478 n984__chipdriverout vss 253.727e-18
c4479 n985__chipdriverout vss 250.42e-18
c4480 n988__chipdriverout vss 175.656e-18
c4481 n989__chipdriverout vss 199.498e-18
c4482 n992__chipdriverout vss 177.656e-18
c4483 n993__chipdriverout vss 218.583e-18
c4484 n996__chipdriverout vss 171.944e-18
c4485 n997__chipdriverout vss 219.459e-18
c4486 n1000__chipdriverout vss 229.173e-18
c4487 n453__i1__i14__net1 vss 38.7349e-18
c4488 n454__i1__i14__net1 vss 34.5754e-18
c4489 n12__i5__i7__y3out vss 115.509e-18
c4490 n13__i5__i7__y0out vss 190.839e-18
c4491 n546__vddio vss 261.328e-18
c4492 n547__vddio vss 259.901e-18
c4493 n550__vddio vss 137.28e-18
c4494 n551__vddio vss 247.956e-18
c4495 n554__vddio vss 142.686e-18
c4496 n555__vddio vss 258.45e-18
c4497 n558__vddio vss 141.176e-18
c4498 n565__vddio vss 193.28e-18
c4499 n939__chipdriverout vss 144.869e-18
c4500 n940__chipdriverout vss 208.199e-18
c4501 n942__chipdriverout vss 176.099e-18
c4502 n943__chipdriverout vss 213.212e-18
c4503 n945__chipdriverout vss 254.179e-18
c4504 n948__chipdriverout vss 245.298e-18
c4505 n951__chipdriverout vss 171.734e-18
c4506 n952__chipdriverout vss 194.419e-18
c4507 n954__chipdriverout vss 173.51e-18
c4508 n955__chipdriverout vss 213.745e-18
c4509 n957__chipdriverout vss 168.068e-18
c4510 n958__chipdriverout vss 214.23e-18
c4511 n960__chipdriverout vss 221.673e-18
c4512 n437__i1__i14__net1 vss 38.6662e-18
c4513 n438__i1__i14__net1 vss 32.9966e-18
c4514 n525__vddio vss 256.719e-18
c4515 n528__vddio vss 253.646e-18
c4516 n529__vddio vss 133.89e-18
c4517 n531__vddio vss 241.726e-18
c4518 n532__vddio vss 139.108e-18
c4519 n534__vddio vss 251.787e-18
c4520 n535__vddio vss 136.945e-18
c4521 n537__vddio vss 160.316e-18
c4522 n900__chipdriverout vss 152.407e-18
c4523 n901__chipdriverout vss 219.247e-18
c4524 n903__chipdriverout vss 183.026e-18
c4525 n904__chipdriverout vss 222.801e-18
c4526 n906__chipdriverout vss 253.738e-18
c4527 n909__chipdriverout vss 257.106e-18
c4528 n912__chipdriverout vss 182.317e-18
c4529 n913__chipdriverout vss 206.705e-18
c4530 n915__chipdriverout vss 183.982e-18
c4531 n916__chipdriverout vss 226.607e-18
c4532 n918__chipdriverout vss 178.086e-18
c4533 n919__chipdriverout vss 225.153e-18
c4534 n921__chipdriverout vss 229.699e-18
c4535 n417__i1__i14__net1 vss 38.7075e-18
c4536 n418__i1__i14__net1 vss 34.3789e-18
c4537 n6__i5__i7__xor2 vss 64.2836e-18
c4538 n8__i5__i7__xor2 vss 77.8475e-18
c4539 n6__i5__i7__xor1 vss 57.2134e-18
c4540 n8__i5__i7__xor1 vss 78.8694e-18
c4541 n504__vddio vss 256.053e-18
c4542 n507__vddio vss 237.935e-18
c4543 n508__vddio vss 134.58e-18
c4544 n510__vddio vss 242.44e-18
c4545 n511__vddio vss 139.678e-18
c4546 n513__vddio vss 251.8e-18
c4547 n514__vddio vss 137.549e-18
c4548 n516__vddio vss 181.913e-18
c4549 n409__i1__i14__net1 vss 43.211e-18
c4550 n410__i1__i14__net1 vss 39.5702e-18
c4551 n884__chipdriverout vss 144.228e-18
c4552 n885__chipdriverout vss 224.253e-18
c4553 n887__chipdriverout vss 192.999e-18
c4554 n888__chipdriverout vss 231.441e-18
c4555 n890__chipdriverout vss 272.825e-18
c4556 n13__i5__i7__x2out vss 114.51e-18
c4557 n13__i5__i7__x1out vss 120.27e-18
c4558 n859__chipdriverout vss 263.602e-18
c4559 n862__chipdriverout vss 204.308e-18
c4560 n863__chipdriverout vss 231.222e-18
c4561 n865__chipdriverout vss 206.594e-18
c4562 n866__chipdriverout vss 218.218e-18
c4563 n868__chipdriverout vss 200.017e-18
c4564 n869__chipdriverout vss 234.744e-18
c4565 n871__chipdriverout vss 263.089e-18
c4566 n16__i5__i7__y2out vss 217.841e-18
c4567 n16__i5__i7__y1out vss 177.105e-18
c4568 n401__i1__i14__net1 vss 46.461e-18
c4569 n402__i1__i14__net1 vss 25.6262e-18
c4570 n483__vddio vss 280.764e-18
c4571 n486__vddio vss 248.593e-18
c4572 n487__vddio vss 155.89e-18
c4573 n489__vddio vss 268.919e-18
c4574 n490__vddio vss 161.629e-18
c4575 n492__vddio vss 247.21e-18
c4576 n493__vddio vss 159.849e-18
c4577 n495__vddio vss 169.16e-18
c4578 n822__chipdriverout vss 149.596e-18
c4579 n823__chipdriverout vss 211.82e-18
c4580 n825__chipdriverout vss 178.239e-18
c4581 n826__chipdriverout vss 216.73e-18
c4582 n828__chipdriverout vss 254.3e-18
c4583 n831__chipdriverout vss 249.075e-18
c4584 n834__chipdriverout vss 175.792e-18
c4585 n835__chipdriverout vss 199.078e-18
c4586 n837__chipdriverout vss 177.638e-18
c4587 n838__chipdriverout vss 218.377e-18
c4588 n840__chipdriverout vss 172.08e-18
c4589 n841__chipdriverout vss 218.966e-18
c4590 n843__chipdriverout vss 225.934e-18
c4591 n14__i5__i7__y2out vss 202.271e-18
c4592 n13__i5__i7__y1out vss 142.744e-18
c4593 n385__i1__i14__net1 vss 46.4771e-18
c4594 n386__i1__i14__net1 vss 23.3097e-18
c4595 n462__vddio vss 272.671e-18
c4596 n465__vddio vss 241.62e-18
c4597 n466__vddio vss 152.13e-18
c4598 n468__vddio vss 262.076e-18
c4599 n469__vddio vss 157.629e-18
c4600 n471__vddio vss 240.168e-18
c4601 n472__vddio vss 156.011e-18
c4602 n474__vddio vss 164.685e-18
c4603 n377__i1__i14__net1 vss 29.79e-18
c4604 n378__i1__i14__net1 vss 40.0651e-18
c4605 n7__i5__i7__y3out vss 110.892e-18
c4606 n5__i5__i7__x3out vss 95.0628e-18
c4607 n783__chipdriverout vss 144.494e-18
c4608 n784__chipdriverout vss 204.652e-18
c4609 n786__chipdriverout vss 172.698e-18
c4610 n787__chipdriverout vss 209.802e-18
c4611 n789__chipdriverout vss 246.277e-18
c4612 n792__chipdriverout vss 249.108e-18
c4613 n795__chipdriverout vss 175.693e-18
c4614 n796__chipdriverout vss 198.951e-18
c4615 n798__chipdriverout vss 177.524e-18
c4616 n799__chipdriverout vss 218.328e-18
c4617 n801__chipdriverout vss 172.055e-18
c4618 n802__chipdriverout vss 219.366e-18
c4619 n804__chipdriverout vss 226.961e-18
c4620 n369__i1__i14__net1 vss 36.3192e-18
c4621 n370__i1__i14__net1 vss 35.8838e-18
c4622 n35__reset vss 45.4322e-18
c4623 n32__reset vss 47.7261e-18
c4624 n435__vddio vss 270.636e-18
c4625 n436__vddio vss 257.684e-18
c4626 n439__vddio vss 136.212e-18
c4627 n440__vddio vss 245.804e-18
c4628 n443__vddio vss 141.492e-18
c4629 n444__vddio vss 256.233e-18
c4630 n447__vddio vss 140.109e-18
c4631 n454__vddio vss 164.58e-18
c4632 n365__i1__i14__net1 vss 43.9303e-18
c4633 n366__i1__i14__net1 vss 49.2928e-18
c4634 n760__chipdriverout vss 220.161e-18
c4635 n762__chipdriverout vss 188.475e-18
c4636 n763__chipdriverout vss 225.429e-18
c4637 n765__chipdriverout vss 265.453e-18
c4638 n742__chipdriverout vss 225.472e-18
c4639 n745__chipdriverout vss 189.36e-18
c4640 n746__chipdriverout vss 212.103e-18
c4641 n748__chipdriverout vss 191.118e-18
c4642 n749__chipdriverout vss 199.197e-18
c4643 n751__chipdriverout vss 185.648e-18
c4644 n752__chipdriverout vss 199.046e-18
c4645 n754__chipdriverout vss 238.74e-18
c4646 n32__i5__i7__i1__net1 vss 195.858e-18
c4647 n75__i5__clk4 vss 99.5439e-18
c4648 n32__i5__i7__i0__net1 vss 134.142e-18
c4649 n74__i5__clk4 vss 96.0239e-18
c4650 n353__i1__i14__net1 vss 28.8673e-18
c4651 n354__i1__i14__net1 vss 35.8995e-18
c4652 n409__vddio vss 283.254e-18
c4653 n412__vddio vss 236.459e-18
c4654 n413__vddio vss 150.363e-18
c4655 n416__vddio vss 257.517e-18
c4656 n417__vddio vss 155.439e-18
c4657 n420__vddio vss 235.008e-18
c4658 n421__vddio vss 154.043e-18
c4659 n433__vddio vss 185.542e-18
c4660 n349__i1__i14__net1 vss 38.9657e-18
c4661 n350__i1__i14__net1 vss 47.238e-18
c4662 n720__chipdriverout vss 149.892e-18
c4663 n721__chipdriverout vss 217.214e-18
c4664 n723__chipdriverout vss 183.039e-18
c4665 n724__chipdriverout vss 222.571e-18
c4666 n726__chipdriverout vss 259.005e-18
c4667 n703__chipdriverout vss 251.456e-18
c4668 n706__chipdriverout vss 178.711e-18
c4669 n707__chipdriverout vss 202.867e-18
c4670 n709__chipdriverout vss 180.689e-18
c4671 n710__chipdriverout vss 222.177e-18
c4672 n712__chipdriverout vss 175.007e-18
c4673 n713__chipdriverout vss 222.459e-18
c4674 n715__chipdriverout vss 231.027e-18
c4675 n337__i1__i14__net1 vss 37.5049e-18
c4676 n338__i1__i14__net1 vss 48.1098e-18
c4677 n59__vdd vss 215.879e-18
c4678 n388__vddio vss 286.555e-18
c4679 n391__vddio vss 240.311e-18
c4680 n392__vddio vss 152.264e-18
c4681 n395__vddio vss 260.735e-18
c4682 n396__vddio vss 157.589e-18
c4683 n399__vddio vss 239.381e-18
c4684 n400__vddio vss 155.318e-18
c4685 n408__vddio vss 164.773e-18
c4686 n329__i1__i14__net1 vss 46.49e-18
c4687 n330__i1__i14__net1 vss 38.6591e-18
c4688 n681__chipdriverout vss 142.918e-18
c4689 n682__chipdriverout vss 199.035e-18
c4690 n684__chipdriverout vss 168.361e-18
c4691 n685__chipdriverout vss 203.997e-18
c4692 n687__chipdriverout vss 241.22e-18
c4693 n664__chipdriverout vss 256.777e-18
c4694 n667__chipdriverout vss 183.389e-18
c4695 n668__chipdriverout vss 208.869e-18
c4696 n670__chipdriverout vss 185.315e-18
c4697 n671__chipdriverout vss 228.248e-18
c4698 n673__chipdriverout vss 179.358e-18
c4699 n674__chipdriverout vss 227.771e-18
c4700 n676__chipdriverout vss 235.109e-18
c4701 n321__i1__i14__net1 vss 22.0834e-18
c4702 n322__i1__i14__net1 vss 46.2093e-18
c4703 n368__vddio vss 265.85e-18
c4704 n369__vddio vss 251.819e-18
c4705 n372__vddio vss 133.724e-18
c4706 n373__vddio vss 239.632e-18
c4707 n376__vddio vss 138.706e-18
c4708 n377__vddio vss 250.972e-18
c4709 n380__vddio vss 137.652e-18
c4710 n387__vddio vss 188.81e-18
c4711 n6__y3 vss 82.3625e-18
c4712 n6__x3 vss 82.8422e-18
c4713 n642__chipdriverout vss 150.703e-18
c4714 n643__chipdriverout vss 212.982e-18
c4715 n645__chipdriverout vss 195.878e-18
c4716 n646__chipdriverout vss 234.399e-18
c4717 n648__chipdriverout vss 253.755e-18
c4718 n625__chipdriverout vss 253.594e-18
c4719 n628__chipdriverout vss 196.565e-18
c4720 n629__chipdriverout vss 222.476e-18
c4721 n631__chipdriverout vss 182.822e-18
c4722 n632__chipdriverout vss 225.442e-18
c4723 n634__chipdriverout vss 176.761e-18
c4724 n635__chipdriverout vss 226.019e-18
c4725 n637__chipdriverout vss 229.741e-18
c4726 n1583__vddio vss 7.14745e-18
c4727 n5__i5__i7__y2out vss 109.583e-18
c4728 n309__i1__i14__net1 vss 24.3913e-18
c4729 n310__i1__i14__net1 vss 31.3084e-18
c4730 n5__i5__i7__x2out vss 101.116e-18
c4731 n347__vddio vss 255.013e-18
c4732 n348__vddio vss 254.928e-18
c4733 n351__vddio vss 134.707e-18
c4734 n352__vddio vss 242.981e-18
c4735 n355__vddio vss 139.933e-18
c4736 n356__vddio vss 253.436e-18
c4737 n359__vddio vss 138.568e-18
c4738 n366__vddio vss 161.737e-18
c4739 n31__reset vss 45.3928e-18
c4740 n29__reset vss 48.3611e-18
c4741 n603__chipdriverout vss 130.883e-18
c4742 n604__chipdriverout vss 227.612e-18
c4743 n606__chipdriverout vss 195.323e-18
c4744 n607__chipdriverout vss 232.951e-18
c4745 n609__chipdriverout vss 271.934e-18
c4746 n586__chipdriverout vss 227.022e-18
c4747 n589__chipdriverout vss 190.418e-18
c4748 n590__chipdriverout vss 214.247e-18
c4749 n592__chipdriverout vss 192.501e-18
c4750 n593__chipdriverout vss 201.138e-18
c4751 n595__chipdriverout vss 186.706e-18
c4752 n596__chipdriverout vss 201.59e-18
c4753 n598__chipdriverout vss 243.012e-18
c4754 n289__i1__i14__net1 vss 24.3913e-18
c4755 n290__i1__i14__net1 vss 32.731e-18
c4756 n28__i5__i7__i1__net1 vss 185.125e-18
c4757 n61__i5__clk4 vss 102.993e-18
c4758 n28__i5__i7__i0__net1 vss 171.173e-18
c4759 n60__i5__clk4 vss 102.938e-18
c4760 n326__vddio vss 274.711e-18
c4761 n329__vddio vss 240.709e-18
c4762 n330__vddio vss 151.804e-18
c4763 n332__vddio vss 261.267e-18
c4764 n333__vddio vss 157.218e-18
c4765 n335__vddio vss 239.258e-18
c4766 n336__vddio vss 155.701e-18
c4767 n338__vddio vss 187.022e-18
c4768 n281__i1__i14__net1 vss 46.4184e-18
c4769 n282__i1__i14__net1 vss 39.755e-18
c4770 n546__chipdriverout vss 131.016e-18
c4771 n549__chipdriverout vss 229.952e-18
c4772 n550__chipdriverout vss 195.74e-18
c4773 n553__chipdriverout vss 234.903e-18
c4774 n554__chipdriverout vss 272.176e-18
c4775 n557__chipdriverout vss 230.255e-18
c4776 n558__chipdriverout vss 193.014e-18
c4777 n561__chipdriverout vss 216.945e-18
c4778 n562__chipdriverout vss 195.008e-18
c4779 n565__chipdriverout vss 203.995e-18
c4780 n566__chipdriverout vss 189.252e-18
c4781 n569__chipdriverout vss 204.254e-18
c4782 n570__chipdriverout vss 245.154e-18
c4783 n61__vdd vss 149.584e-18
c4784 n305__vddio vss 265.813e-18
c4785 n306__vddio vss 253.929e-18
c4786 n309__vddio vss 135.016e-18
c4787 n310__vddio vss 241.917e-18
c4788 n313__vddio vss 139.984e-18
c4789 n314__vddio vss 253.124e-18
c4790 n317__vddio vss 139.029e-18
c4791 n324__vddio vss 164.524e-18
c4792 n265__i1__i14__net1 vss 46.4184e-18
c4793 n266__i1__i14__net1 vss 47.2502e-18
c4794 n59__i5__clk4 vss 437.213e-18
c4795 n27__i5__i7__i1__net1 vss 175.152e-18
c4796 n58__i5__clk4 vss 423.275e-18
c4797 n510__chipdriverout vss 228.795e-18
c4798 n511__chipdriverout vss 195.762e-18
c4799 n514__chipdriverout vss 234.264e-18
c4800 n515__chipdriverout vss 272.196e-18
c4801 n518__chipdriverout vss 233.971e-18
c4802 n519__chipdriverout vss 199.107e-18
c4803 n522__chipdriverout vss 224.99e-18
c4804 n523__chipdriverout vss 201.228e-18
c4805 n526__chipdriverout vss 212.119e-18
c4806 n527__chipdriverout vss 195.009e-18
c4807 n530__chipdriverout vss 212.297e-18
c4808 n531__chipdriverout vss 251.539e-18
c4809 n261__i1__i14__net1 vss 30.7112e-18
c4810 n262__i1__i14__net1 vss 37.302e-18
c4811 n284__vddio vss 263.398e-18
c4812 n287__vddio vss 251.634e-18
c4813 n288__vddio vss 133.625e-18
c4814 n290__vddio vss 239.431e-18
c4815 n291__vddio vss 138.591e-18
c4816 n293__vddio vss 250.565e-18
c4817 n294__vddio vss 137.524e-18
c4818 n296__vddio vss 188.218e-18
c4819 n6__y2 vss 89.2968e-18
c4820 n6__x2 vss 86.7378e-18
c4821 n486__chipdriverout vss 131.649e-18
c4822 n487__chipdriverout vss 231.096e-18
c4823 n489__chipdriverout vss 197.649e-18
c4824 n490__chipdriverout vss 236.554e-18
c4825 n492__chipdriverout vss 276.472e-18
c4826 n469__chipdriverout vss 233.593e-18
c4827 n472__chipdriverout vss 198.24e-18
c4828 n473__chipdriverout vss 223.652e-18
c4829 n475__chipdriverout vss 200.254e-18
c4830 n476__chipdriverout vss 210.875e-18
c4831 n478__chipdriverout vss 193.667e-18
c4832 n479__chipdriverout vss 209.845e-18
c4833 n481__chipdriverout vss 250.868e-18
c4834 n245__i1__i14__net1 vss 30.512e-18
c4835 n246__i1__i14__net1 vss 37.3412e-18
c4836 n2__i5__i7__y1out vss 69.5796e-18
c4837 n2__i5__i7__x1out vss 64.5725e-18
c4838 n253__vddio vss 277.994e-18
c4839 n256__vddio vss 232.141e-18
c4840 n257__vddio vss 147.971e-18
c4841 n259__vddio vss 252.554e-18
c4842 n260__vddio vss 153.019e-18
c4843 n262__vddio vss 231.102e-18
c4844 n263__vddio vss 150.893e-18
c4845 n265__vddio vss 179.435e-18
c4846 n233__i1__i14__net1 vss 38.4703e-18
c4847 n234__i1__i14__net1 vss 37.4507e-18
c4848 n21__reset vss 45.6881e-18
c4849 n20__reset vss 47.0051e-18
c4850 n432__chipdriverout vss 131.04e-18
c4851 n433__chipdriverout vss 221.37e-18
c4852 n435__chipdriverout vss 190.223e-18
c4853 n436__chipdriverout vss 226.812e-18
c4854 n438__chipdriverout vss 261.384e-18
c4855 n441__chipdriverout vss 229.809e-18
c4856 n444__chipdriverout vss 196.803e-18
c4857 n445__chipdriverout vss 221.905e-18
c4858 n447__chipdriverout vss 199.142e-18
c4859 n448__chipdriverout vss 208.484e-18
c4860 n450__chipdriverout vss 193.066e-18
c4861 n451__chipdriverout vss 210.476e-18
c4862 n453__chipdriverout vss 252.447e-18
c4863 n229__i1__i14__net1 vss 30.4688e-18
c4864 n230__i1__i14__net1 vss 40.0859e-18
c4865 n232__vddio vss 274.873e-18
c4866 n233__vddio vss 262.482e-18
c4867 n236__vddio vss 138.516e-18
c4868 n237__vddio vss 250.45e-18
c4869 n240__vddio vss 144.073e-18
c4870 n241__vddio vss 261.031e-18
c4871 n244__vddio vss 142.413e-18
c4872 n251__vddio vss 166.95e-18
c4873 n23__i5__i7__i1__net1 vss 184.96e-18
c4874 n52__i5__clk4 vss 104.473e-18
c4875 n23__i5__i7__i0__net1 vss 169.392e-18
c4876 n50__i5__clk4 vss 108.439e-18
c4877 n221__i1__i14__net1 vss 46.6327e-18
c4878 n222__i1__i14__net1 vss 37.2498e-18
c4879 n393__chipdriverout vss 128.487e-18
c4880 n394__chipdriverout vss 219.394e-18
c4881 n396__chipdriverout vss 188.71e-18
c4882 n397__chipdriverout vss 224.487e-18
c4883 n399__chipdriverout vss 263.409e-18
c4884 n402__chipdriverout vss 224.307e-18
c4885 n405__chipdriverout vss 189.611e-18
c4886 n406__chipdriverout vss 213.337e-18
c4887 n408__chipdriverout vss 191.664e-18
c4888 n409__chipdriverout vss 200.359e-18
c4889 n411__chipdriverout vss 185.899e-18
c4890 n412__chipdriverout vss 200.75e-18
c4891 n414__chipdriverout vss 240.85e-18
c4892 n213__i1__i14__net1 vss 29.3252e-18
c4893 n214__i1__i14__net1 vss 38.6834e-18
c4894 n211__vddio vss 283.699e-18
c4895 n214__vddio vss 237.097e-18
c4896 n215__vddio vss 149.506e-18
c4897 n217__vddio vss 257.411e-18
c4898 n218__vddio vss 154.912e-18
c4899 n220__vddio vss 235.605e-18
c4900 n221__vddio vss 153.311e-18
c4901 n223__vddio vss 160.604e-18
c4902 n354__chipdriverout vss 144.652e-18
c4903 n355__chipdriverout vss 218.46e-18
c4904 n357__chipdriverout vss 188.188e-18
c4905 n358__chipdriverout vss 223.644e-18
c4906 n360__chipdriverout vss 263.237e-18
c4907 n363__chipdriverout vss 231.528e-18
c4908 n366__chipdriverout vss 196.522e-18
c4909 n367__chipdriverout vss 222.116e-18
c4910 n369__chipdriverout vss 198.672e-18
c4911 n370__chipdriverout vss 209.118e-18
c4912 n372__chipdriverout vss 192.469e-18
c4913 n373__chipdriverout vss 209.347e-18
c4914 n375__chipdriverout vss 248.181e-18
c4915 n45__i5__clk4 vss 443.621e-18
c4916 n44__i5__clk4 vss 435.988e-18
c4917 n180__vddio vss 283.823e-18
c4918 n183__vddio vss 234.556e-18
c4919 n184__vddio vss 148.748e-18
c4920 n186__vddio vss 254.755e-18
c4921 n187__vddio vss 153.976e-18
c4922 n189__vddio vss 233.708e-18
c4923 n190__vddio vss 152.631e-18
c4924 n192__vddio vss 160.653e-18
c4925 n189__i1__i14__net1 vss 39.1512e-18
c4926 n190__i1__i14__net1 vss 46.2987e-18
c4927 n315__chipdriverout vss 128.548e-18
c4928 n316__chipdriverout vss 219.534e-18
c4929 n318__chipdriverout vss 188.77e-18
c4930 n319__chipdriverout vss 224.676e-18
c4931 n321__chipdriverout vss 263.29e-18
c4932 n324__chipdriverout vss 235.079e-18
c4933 n327__chipdriverout vss 199.643e-18
c4934 n328__chipdriverout vss 225.246e-18
c4935 n330__chipdriverout vss 201.711e-18
c4936 n331__chipdriverout vss 213.598e-18
c4937 n333__chipdriverout vss 195.743e-18
c4938 n334__chipdriverout vss 213.315e-18
c4939 n336__chipdriverout vss 256.415e-18
c4940 n7__y1 vss 81.294e-18
c4941 n6__x1 vss 81.2927e-18
c4942 n1591__vddio vss 7.44695e-18
c4943 n181__i1__i14__net1 vss 31.104e-18
c4944 n182__i1__i14__net1 vss 26.125e-18
c4945 n159__vddio vss 271.284e-18
c4946 n162__vddio vss 237.198e-18
c4947 n163__vddio vss 134.625e-18
c4948 n165__vddio vss 241.179e-18
c4949 n166__vddio vss 155.39e-18
c4950 n168__vddio vss 236.268e-18
c4951 n169__vddio vss 153.96e-18
c4952 n171__vddio vss 185.961e-18
c4953 n2__i5__i7__y0out vss 104.809e-18
c4954 n2__i5__i7__x0out vss 99.463e-18
c4955 n276__chipdriverout vss 16.859e-18
c4956 n277__chipdriverout vss 203.255e-18
c4957 n279__chipdriverout vss 188.771e-18
c4958 n280__chipdriverout vss 224.424e-18
c4959 n282__chipdriverout vss 246.779e-18
c4960 n285__chipdriverout vss 250.862e-18
c4961 n288__chipdriverout vss 192.759e-18
c4962 n289__chipdriverout vss 216.587e-18
c4963 n291__chipdriverout vss 178.619e-18
c4964 n292__chipdriverout vss 219.133e-18
c4965 n294__chipdriverout vss 173.106e-18
c4966 n295__chipdriverout vss 219.163e-18
c4967 n297__chipdriverout vss 228.09e-18
c4968 n165__i1__i14__net1 vss 24.8261e-18
c4969 n166__i1__i14__net1 vss 47.1219e-18
c4970 n12__reset vss 45.5815e-18
c4971 n9__reset vss 46.805e-18
c4972 n138__vddio vss 268.442e-18
c4973 n141__vddio vss 255.922e-18
c4974 n142__vddio vss 135.416e-18
c4975 n144__vddio vss 243.56e-18
c4976 n145__vddio vss 139.965e-18
c4977 n147__vddio vss 253.812e-18
c4978 n148__vddio vss 138.515e-18
c4979 n150__vddio vss 162.64e-18
c4980 n153__i1__i14__net1 vss 39.1009e-18
c4981 n154__i1__i14__net1 vss 46.0657e-18
c4982 n14__i5__i7__i1__net1 vss 183.959e-18
c4983 n33__i5__clk4 vss 91.2077e-18
c4984 n14__i5__i7__i0__net1 vss 161.502e-18
c4985 n32__i5__clk4 vss 96.1353e-18
c4986 n237__chipdriverout vss 145.515e-18
c4987 n238__chipdriverout vss 203.255e-18
c4988 n240__chipdriverout vss 172.399e-18
c4989 n241__chipdriverout vss 208.283e-18
c4990 n243__chipdriverout vss 246.779e-18
c4991 n246__chipdriverout vss 247.083e-18
c4992 n249__chipdriverout vss 173.888e-18
c4993 n250__chipdriverout vss 197.175e-18
c4994 n252__chipdriverout vss 175.734e-18
c4995 n253__chipdriverout vss 215.695e-18
c4996 n255__chipdriverout vss 170.191e-18
c4997 n256__chipdriverout vss 216.514e-18
c4998 n258__chipdriverout vss 224.863e-18
c4999 n149__i1__i14__net1 vss 24.8261e-18
c5000 n150__i1__i14__net1 vss 47.1219e-18
c5001 n65__vdd vss 191.841e-18
c5002 n117__vddio vss 265.75e-18
c5003 n120__vddio vss 253.067e-18
c5004 n121__vddio vss 133.654e-18
c5005 n123__vddio vss 240.561e-18
c5006 n124__vddio vss 138.188e-18
c5007 n126__vddio vss 251.575e-18
c5008 n127__vddio vss 136.821e-18
c5009 n129__vddio vss 182.778e-18
c5010 n137__i1__i14__net1 vss 44.8806e-18
c5011 n138__i1__i14__net1 vss 35.7489e-18
c5012 n198__chipdriverout vss 151.553e-18
c5013 n199__chipdriverout vss 215.829e-18
c5014 n201__chipdriverout vss 182.574e-18
c5015 n202__chipdriverout vss 221.033e-18
c5016 n204__chipdriverout vss 258.19e-18
c5017 n207__chipdriverout vss 248.606e-18
c5018 n210__chipdriverout vss 175.962e-18
c5019 n211__chipdriverout vss 201.099e-18
c5020 n213__chipdriverout vss 178.048e-18
c5021 n214__chipdriverout vss 218.669e-18
c5022 n216__chipdriverout vss 171.735e-18
c5023 n217__chipdriverout vss 219.995e-18
c5024 n219__chipdriverout vss 226.966e-18
c5025 n129__i1__i14__net1 vss 25.9367e-18
c5026 n130__i1__i14__net1 vss 34.2481e-18
c5027 n96__vddio vss 255.205e-18
c5028 n99__vddio vss 252.692e-18
c5029 n100__vddio vss 133.868e-18
c5030 n102__vddio vss 240.291e-18
c5031 n103__vddio vss 138.161e-18
c5032 n105__vddio vss 251.128e-18
c5033 n106__vddio vss 137.077e-18
c5034 n108__vddio vss 161.141e-18
c5035 n31__i5__clk4 vss 345.317e-18
c5036 n13__i5__i7__i1__net1 vss 164.882e-18
c5037 n30__i5__clk4 vss 255.772e-18
c5038 n159__chipdriverout vss 151.203e-18
c5039 n160__chipdriverout vss 212.322e-18
c5040 n162__chipdriverout vss 179.324e-18
c5041 n163__chipdriverout vss 217.52e-18
c5042 n165__chipdriverout vss 255.862e-18
c5043 n168__chipdriverout vss 262.579e-18
c5044 n171__chipdriverout vss 185.97e-18
c5045 n172__chipdriverout vss 211.141e-18
c5046 n174__chipdriverout vss 187.751e-18
c5047 n175__chipdriverout vss 229.665e-18
c5048 n177__chipdriverout vss 181.838e-18
c5049 n178__chipdriverout vss 230.637e-18
c5050 n180__chipdriverout vss 237.507e-18
c5051 n117__i1__i14__net1 vss 33.2171e-18
c5052 n118__i1__i14__net1 vss 27.34e-18
c5053 n6__y0 vss 79.73e-18
c5054 n6__x0 vss 81.6023e-18
c5055 n69__vddio vss 283.24e-18
c5056 n72__vddio vss 248.593e-18
c5057 n73__vddio vss 155.951e-18
c5058 n75__vddio vss 268.367e-18
c5059 n76__vddio vss 161.087e-18
c5060 n78__vddio vss 247.21e-18
c5061 n79__vddio vss 159.308e-18
c5062 n81__vddio vss 191.74e-18
c5063 n109__i1__i14__net1 vss 36.4148e-18
c5064 n110__i1__i14__net1 vss 48.8694e-18
c5065 n135__chipdriverout vss 134.796e-18
c5066 n136__chipdriverout vss 228.696e-18
c5067 n138__chipdriverout vss 196.136e-18
c5068 n139__chipdriverout vss 234.114e-18
c5069 n141__chipdriverout vss 273.071e-18
c5070 n118__chipdriverout vss 226.21e-18
c5071 n121__chipdriverout vss 191.664e-18
c5072 n122__chipdriverout vss 215.39e-18
c5073 n124__chipdriverout vss 193.718e-18
c5074 n125__chipdriverout vss 201.571e-18
c5075 n127__chipdriverout vss 188.031e-18
c5076 n128__chipdriverout vss 202.324e-18
c5077 n130__chipdriverout vss 243.5e-18
c5078 n7__i5__i7__i1__net1 vss 53.4265e-18
c5079 n7__i5__i7__i0__net1 vss 37.9827e-18
c5080 n101__i1__i14__net1 vss 32.2596e-18
c5081 n102__i1__i14__net1 vss 24.9976e-18
c5082 n23__i5__clk4 vss 197.989e-18
c5083 n22__i5__clk4 vss 226.748e-18
c5084 n44__vddio vss 278.869e-18
c5085 n47__vddio vss 241.62e-18
c5086 n48__vddio vss 152.13e-18
c5087 n50__vddio vss 261.436e-18
c5088 n51__vddio vss 156.994e-18
c5089 n53__vddio vss 240.168e-18
c5090 n54__vddio vss 155.376e-18
c5091 n56__vddio vss 187.157e-18
c5092 n93__i1__i14__net1 vss 43.5539e-18
c5093 n94__i1__i14__net1 vss 39.8464e-18
c5094 n96__chipdriverout vss 134.642e-18
c5095 n97__chipdriverout vss 228.055e-18
c5096 n99__chipdriverout vss 195.608e-18
c5097 n100__chipdriverout vss 233.434e-18
c5098 n102__chipdriverout vss 272.839e-18
c5099 n79__chipdriverout vss 226.198e-18
c5100 n82__chipdriverout vss 191.725e-18
c5101 n83__chipdriverout vss 215.451e-18
c5102 n85__chipdriverout vss 193.779e-18
c5103 n86__chipdriverout vss 201.571e-18
c5104 n88__chipdriverout vss 188.091e-18
c5105 n89__chipdriverout vss 202.324e-18
c5106 n91__chipdriverout vss 243.727e-18
c5107 n23__vddio vss 278.65e-18
c5108 n26__vddio vss 241.491e-18
c5109 n27__vddio vss 152.13e-18
c5110 n29__vddio vss 261.343e-18
c5111 n30__vddio vss 156.868e-18
c5112 n32__vddio vss 240.014e-18
c5113 n33__vddio vss 154.969e-18
c5114 n35__vddio vss 164.144e-18
c5115 n73__i1__i14__net1 vss 36.3698e-18
c5116 n74__i1__i14__net1 vss 48.6706e-18
c5117 n58__chipdriverout vss 229.279e-18
c5118 n60__chipdriverout vss 196.78e-18
c5119 n61__chipdriverout vss 234.643e-18
c5120 n63__chipdriverout vss 273.227e-18
c5121 n40__chipdriverout vss 226.438e-18
c5122 n43__chipdriverout vss 192.2e-18
c5123 n44__chipdriverout vss 216.041e-18
c5124 n46__chipdriverout vss 194.263e-18
c5125 n47__chipdriverout vss 202.122e-18
c5126 n49__chipdriverout vss 188.235e-18
c5127 n50__chipdriverout vss 202.742e-18
c5128 n52__chipdriverout vss 242.668e-18
c5129 n69__i1__i14__net1 vss 34.2388e-18
c5130 n70__i1__i14__net1 vss 26.7035e-18
c5131 n2__vddio vss 274.514e-18
c5132 n5__vddio vss 241.099e-18
c5133 n6__vddio vss 156.513e-18
c5134 n8__vddio vss 265.674e-18
c5135 n9__vddio vss 161.264e-18
c5136 n11__vddio vss 239.227e-18
c5137 n12__vddio vss 159.017e-18
c5138 n14__vddio vss 235.347e-18
c5139 n62__i1__i14__net1 vss 48.08e-18
c5140 n61__i1__i14__net1 vss 33.4575e-18
c5141 n18__chipdriverout vss 91.3774e-18
c5142 n19__chipdriverout vss 154.193e-18
c5143 n21__chipdriverout vss 130.469e-18
c5144 n22__chipdriverout vss 157.022e-18
c5145 n24__chipdriverout vss 183.943e-18
c5146 n14__chipdriverout vss 166.408e-18
c5147 n12__chipdriverout vss 136.469e-18
c5148 n11__chipdriverout vss 153.573e-18
c5149 n9__chipdriverout vss 137.162e-18
c5150 n8__chipdriverout vss 148.138e-18
c5151 n6__chipdriverout vss 134.233e-18
c5152 n5__chipdriverout vss 149.099e-18
c5153 n2__chipdriverout vss 175.075e-18
c5154 n1631__vddio vss 33.3158e-15
c5155 n1767__vddio vss 655.336e-18
c5156 n1815__vddio vss 114.073e-18
c5157 n187__i1__i13__net1 vss 340.489e-18
c5158 n1807__vddio vss 227.097e-18
c5159 n176__i1__i13__net1 vss 336.815e-18
c5160 n1800__vddio vss 226.149e-18
c5161 n165__i1__i13__net1 vss 344.535e-18
c5162 n1794__vddio vss 131.529e-18
c5163 n1786__vddio vss 109.08e-18
c5164 n1766__vddio vss 55.7464e-18
c5165 n326__i1__net2 vss 306.731e-18
c5166 n26__i1__net4 vss 177.13e-18
c5167 n1760__vddio vss 223.517e-18
c5168 n1776__vddio vss 55.6366e-18
c5169 n317__i1__net2 vss 302.511e-18
c5170 n1753__vddio vss 222.244e-18
c5171 n304__i1__net2 vss 309.943e-18
c5172 n1784__vddio vss 56.6968e-18
c5173 n1746__vddio vss 228.439e-18
c5174 n8__i1__i11__outinv vss 175.128e-18
c5175 n295__i1__net2 vss 322.922e-18
c5176 n1778__vddio vss 81.7886e-18
c5177 n1739__vddio vss 229.843e-18
c5178 n181__i1__i13__net1 vss 236.482e-18
c5179 n170__i1__i13__net1 vss 240.203e-18
c5180 n159__i1__i13__net1 vss 234.415e-18
c5181 n320__i1__net2 vss 214.674e-18
c5182 n27__i1__net4 vss 153.181e-18
c5183 n311__i1__net2 vss 221.691e-18
c5184 n24__i1__net4 vss 126.181e-18
c5185 n307__i1__net2 vss 218.888e-18
c5186 n5__i1__i11__outinv vss 142.389e-18
c5187 n298__i1__net2 vss 244.668e-18
c5188 n9__i1__i11__outinv vss 99.9175e-18
c5189 n289__i1__net2 vss 234.4e-18
c5190 n280__i1__net2 vss 242.201e-18
c5191 n271__i1__net2 vss 239.149e-18
c5192 n29__i1__net3 vss 199.104e-18
c5193 n262__i1__net2 vss 232.24e-18
c5194 n253__i1__net2 vss 233.837e-18
c5195 n9__i1__net3 vss 42.246e-21
c5196 n239__i1__net2 vss 243.131e-18
c5197 n235__i1__net2 vss 140.44e-18
c5198 n286__i1__net2 vss 309.095e-18
c5199 n1779__vddio vss 151.799e-18
c5200 n1714__vddio vss 226.259e-18
c5201 n277__i1__net2 vss 304.091e-18
c5202 n1780__vddio vss 159.89e-18
c5203 n1708__vddio vss 229.754e-18
c5204 n268__i1__net2 vss 309.796e-18
c5205 n1781__vddio vss 154.096e-18
c5206 n1700__vddio vss 226.418e-18
c5207 n259__i1__net2 vss 300.35e-18
c5208 n1782__vddio vss 250.701e-18
c5209 n1693__vddio vss 222.834e-18
c5210 n19__i1__net3 vss 410.471e-24
c5211 n250__i1__net2 vss 306.501e-18
c5212 n1783__vddio vss 256.028e-18
c5213 n1686__vddio vss 227.829e-18
c5214 n12__i1__net3 vss 151.846e-21
c5215 n245__i1__net2 vss 305.408e-18
c5216 n1775__vddio vss 279.87e-18
c5217 n1679__vddio vss 223.96e-18
c5218 n232__i1__net2 vss 184.559e-18
c5219 n1523__vddio vss 244.701e-18
c5220 n44__shift vss 54.9604e-18
c5221 n1331__i1__i14__net1 vss 397.964e-18
c5222 n375__vdd vss 66.6934e-18
c5223 n181__vdd vss 83.0464e-18
c5224 n4__piso_outinv vss 87.7588e-18
c5225 n1487__vddio vss 419.52e-18
c5226 n374__vdd vss 85.9114e-18
c5227 n4__i5__i8__i8__net1 vss 76.9116e-18
c5228 n8__piso_outinv vss 83.4551e-18
c5229 n1272__i1__i14__net1 vss 394.149e-18
c5230 n372__vdd vss 66.4912e-18
c5231 n269__vdd vss 78.6743e-18
c5232 n46__shift vss 32.8953e-18
c5233 n182__vdd vss 1.39376e-15
c5234 n1325__i1__i14__net1 vss 285.615e-18
c5235 n328__vdd vss 2.35719e-15
c5236 n7__piso_outinv vss 55.3455e-18
c5237 n6__piso_outinv vss 45.6102e-18
c5238 n1260__i1__i14__net1 vss 284.303e-18
c5239 n6__i5__i8__i8__net1 vss 54.2238e-18
c5240 n1453__vddio vss 408.594e-18
c5241 n370__vdd vss 58.439e-18
c5242 n1222__i1__i14__net1 vss 371.61e-18
c5243 n14__piso_out vss 95.8624e-18
c5244 n13__i5__i8__net5 vss 41.3569e-18
c5245 n368__vdd vss 72.6153e-18
c5246 n270__vdd vss 66.3574e-18
c5247 n1432__vddio vss 404.44e-18
c5248 n18__i5__i8__net5 vss 59.5225e-18
c5249 n7__i4__net1 vss 70.9454e-18
c5250 n271__vdd vss 43.7972e-18
c5251 n1183__i1__i14__net1 vss 370.345e-18
c5252 n365__vdd vss 59.3197e-18
c5253 n1236__i1__i14__net1 vss 283.103e-18
c5254 n17__piso_out vss 61.6246e-18
c5255 n17__i5__i8__net5 vss 31.9247e-18
c5256 n16__i5__i8__net5 vss 43.8061e-18
c5257 n9__i4__net1 vss 44.3191e-18
c5258 n1197__i1__i14__net1 vss 283.386e-18
c5259 n95__i5__clk4 vss 61.4337e-18
c5260 n4__bufin vss 64.9228e-18
c5261 n1143__i1__i14__net1 vss 411.311e-18
c5262 n96__i5__clk4 vss 66.9541e-18
c5263 n9__bufin vss 69.2083e-18
c5264 n7__i5__i8__i10__net23 vss 101.449e-21
c5265 n8__i5__i6__i5__net23 vss 29.5554e-21
c5266 n1104__i1__i14__net1 vss 283.31e-18
c5267 n93__i5__clk4 vss 69.0974e-18
c5268 n8__bufin vss 73.2446e-18
c5269 n4__i5__i8__i10__net23 vss 112.077e-21
c5270 n4__i5__i6__i5__net23 vss 242.047e-21
c5271 n1098__i1__i14__net1 vss 283.277e-18
c5272 n8__i5__i8__i10__net21 vss 105.992e-21
c5273 n8__i5__i6__i5__net21 vss 9.1938e-21
c5274 n10__i5__i8__i10__net22 vss 70.0209e-18
c5275 n10__i5__i6__i5__net22 vss 69.6373e-18
c5276 n1041__i1__i14__net1 vss 295.644e-18
c5277 n4__i5__i8__i10__net21 vss 112.077e-21
c5278 n1411__vddio vss 414.159e-18
c5279 n1155__i1__i14__net1 vss 392.315e-18
c5280 n1380__vddio vss 417.896e-18
c5281 n7__i5__i8__i10__net24 vss 40.9775e-18
c5282 n8__i5__i6__i5__net24 vss 39.9707e-18
c5283 n1116__i1__i14__net1 vss 393.993e-18
c5284 n97__i5__clk4 vss 111.097e-18
c5285 n10__bufin vss 113.17e-18
c5286 n4__i5__i8__i10__net24 vss 60.4273e-18
c5287 n4__i5__i6__i5__net24 vss 60.5458e-18
c5288 n1359__vddio vss 408.538e-18
c5289 n272__vdd vss 116.715e-18
c5290 n362__vdd vss 117.328e-18
c5291 n1091__i1__i14__net1 vss 371.61e-18
c5292 n1351__vddio vss 404.44e-18
c5293 n8__i5__i8__i10__net25 vss 48.8267e-18
c5294 n8__i5__i6__i5__net25 vss 45.819e-18
c5295 n8__i5__i8__i10__net22 vss 124.942e-18
c5296 n8__i5__i6__i5__net22 vss 115.369e-18
c5297 n1027__i1__i14__net1 vss 384.652e-18
c5298 n4__i5__i8__i10__net25 vss 61.5921e-18
c5299 n4__i5__i6__i5__net25 vss 63.0529e-18
c5300 n273__vdd vss 123.141e-18
c5301 n359__vdd vss 118.135e-18
c5302 n1317__vddio vss 409.618e-18
c5303 n987__i1__i14__net1 vss 271.965e-18
c5304 n8__i5__i6__net35 vss 34.1859e-18
c5305 n22__i5__i8__net1 vss 31.7369e-18
c5306 n13__i5__r0 vss 60.7086e-18
c5307 n21__i5__i8__net1 vss 42.5959e-18
c5308 n948__i1__i14__net1 vss 406.817e-18
c5309 n14__i5__i6__net35 vss 68.6306e-18
c5310 n10__i5__i6__net34 vss 47.0771e-18
c5311 n999__i1__i14__net1 vss 394.149e-18
c5312 n10__i5__i6__net35 vss 151.092e-18
c5313 n18__i5__i8__net1 vss 46.0137e-18
c5314 n1296__vddio vss 418.026e-18
c5315 n11__i5__r0 vss 70.6287e-18
c5316 n274__vdd vss 69.6165e-18
c5317 n23__i5__i8__net1 vss 59.4174e-18
c5318 n960__i1__i14__net1 vss 392.49e-18
c5319 n12__i5__i6__net35 vss 179.986e-18
c5320 n275__vdd vss 43.6785e-18
c5321 n9__i5__i6__net34 vss 53.2521e-18
c5322 n1265__vddio vss 413.899e-18
c5323 n7__i5__i6__i8__net4 vss 104.718e-18
c5324 n921__i1__i14__net1 vss 388.435e-18
c5325 n356__vdd vss 59.7538e-18
c5326 n26__i5__i8__net2 vss 47.7941e-18
c5327 n5__i5__i6__i8__net4 vss 157.567e-18
c5328 n909__i1__i14__net1 vss 406.79e-18
c5329 n28__i5__i8__net2 vss 69.185e-18
c5330 n870__i1__i14__net1 vss 271.763e-18
c5331 n8__i5__i8__i9__net23 vss 102.312e-21
c5332 n25__i5__i8__net2 vss 72.6697e-18
c5333 n6__i5__i6__net34 vss 71.4988e-18
c5334 n4__i5__i8__i9__net23 vss 112.077e-21
c5335 n831__i1__i14__net1 vss 270.596e-18
c5336 n7__i5__i6__i4__net23 vss 102.844e-21
c5337 n5__i5__i6__net34 vss 74.2932e-18
c5338 n4__i5__i6__i4__net23 vss 90.5897e-21
c5339 n7__i5__i8__i9__net21 vss 106.854e-21
c5340 n792__i1__i14__net1 vss 273.739e-18
c5341 n10__i5__i8__i9__net22 vss 71.0337e-18
c5342 n4__i5__i8__i9__net21 vss 112.077e-21
c5343 n7__i5__i6__i4__net21 vss 124.143e-21
c5344 n1257__vddio vss 405.301e-18
c5345 n882__i1__i14__net1 vss 390.242e-18
c5346 n8__i5__i8__i9__net24 vss 46.1535e-18
c5347 n29__i5__i8__net2 vss 111.682e-18
c5348 n1223__vddio vss 409.66e-18
c5349 n4__i5__i8__i9__net24 vss 60.8347e-18
c5350 n276__vdd vss 117.073e-18
c5351 n843__i1__i14__net1 vss 395.592e-18
c5352 n7__i5__i6__i4__net24 vss 41.0307e-18
c5353 n7__i5__i6__net34 vss 111.997e-18
c5354 n1202__vddio vss 419.48e-18
c5355 n4__i5__i6__i4__net24 vss 60.0367e-18
c5356 n7__i5__i8__i9__net25 vss 46.4613e-18
c5357 n353__vdd vss 117.933e-18
c5358 n804__i1__i14__net1 vss 397.115e-18
c5359 n8__i5__i8__i9__net22 vss 117.37e-18
c5360 n4__i5__i8__i9__net25 vss 62.5531e-18
c5361 n1175__vddio vss 226.799e-18
c5362 n277__vdd vss 116.914e-18
c5363 n7__i5__i6__i4__net25 vss 45.6135e-18
c5364 n8__i5__i6__i4__net22 vss 115.02e-18
c5365 n10__i5__i6__i4__net22 vss 71.6879e-18
c5366 n4__i5__i6__i4__net21 vss 149.084e-21
c5367 n13__i5__i8__net4 vss 42.5056e-18
c5368 n4__i5__i6__i4__net25 vss 62.7037e-18
c5369 n8__i5__i8__net4 vss 46.8811e-18
c5370 n350__vdd vss 118.242e-18
c5371 n278__vdd vss 73.5089e-18
c5372 n14__i5__i8__net4 vss 61.5366e-18
c5373 n11__i5__i8__net4 vss 42.7182e-18
c5374 n8__i5__i6__net33 vss 34.7057e-18
c5375 n279__vdd vss 38.4525e-18
c5376 n10__i5__i6__net33 vss 150.381e-18
c5377 n10__i5__r1 vss 70.553e-18
c5378 n161__vdd vss 27.8816e-18
c5379 n12__i5__i6__net33 vss 178.61e-18
c5380 n49__i5__clk_buf vss 116.027e-18
c5381 n9__i5__i6__net32 vss 53.3085e-18
c5382 n155__vdd vss 68.1623e-18
c5383 n1101__vddio vss 226.871e-18
c5384 n50__i5__clk_buf vss 116.496e-18
c5385 n7__i5__i6__i7__net4 vss 105.297e-18
c5386 n1892__chipdriverout vss 373.193e-18
c5387 n152__vdd vss 125.204e-21
c5388 n347__vdd vss 61.0153e-18
c5389 n12__i5__r1 vss 60.5044e-18
c5390 n14__i5__i6__net33 vss 68.3429e-18
c5391 n48__i5__clk_buf vss 73.6619e-18
c5392 n10__i5__i6__net32 vss 46.7523e-18
c5393 n47__i5__clk_buf vss 72.8535e-18
c5394 n5__i5__i6__i7__net4 vss 156.277e-18
c5395 n1906__chipdriverout vss 417.113e-18
c5396 n20__i5__i9__net21 vss 59.9728e-18
c5397 n1867__chipdriverout vss 291.86e-18
c5398 n6__i5__i6__net32 vss 70.8062e-18
c5399 n1080__vddio vss 405.885e-18
c5400 n280__vdd vss 59.2144e-18
c5401 n18__i5__i9__net21 vss 102.723e-18
c5402 n1853__chipdriverout vss 385.294e-18
c5403 n281__vdd vss 78.4058e-18
c5404 n1059__vddio vss 431.499e-18
c5405 n7__i5__i6__i2__net24 vss 41.1256e-18
c5406 n10__i5__r2 vss 42.3559e-18
c5407 n1830__chipdriverout vss 361.971e-18
c5408 n7__i5__i6__net32 vss 110.076e-18
c5409 n282__vdd vss 58.3616e-18
c5410 n7__i5__i6__i2__net23 vss 1.18871e-18
c5411 n11__i5__r2 vss 51.6272e-18
c5412 n1823__chipdriverout vss 278.603e-18
c5413 n5__i5__i6__net32 vss 76.8605e-18
c5414 n4__i5__i6__i2__net24 vss 60.161e-18
c5415 n1038__vddio vss 412.398e-18
c5416 n344__vdd vss 117.624e-18
c5417 n1775__chipdriverout vss 366.318e-18
c5418 n283__vdd vss 65.0207e-18
c5419 n1020__vddio vss 394.876e-18
c5420 n7__i5__i6__i2__net25 vss 45.6008e-18
c5421 n8__i5__i6__i2__net22 vss 113.659e-18
c5422 n1736__chipdriverout vss 370.634e-18
c5423 n4__i5__i6__i2__net25 vss 62.7597e-18
c5424 n4__i5__i7__i7__net3 vss 319.892e-18
c5425 n986__vddio vss 403.879e-18
c5426 n341__vdd vss 118.388e-18
c5427 n1697__chipdriverout vss 377.895e-18
c5428 n4__i5__i6__i2__net23 vss 1.75157e-18
c5429 n1789__chipdriverout vss 278.505e-18
c5430 n7__i5__i6__i2__net21 vss 727.081e-21
c5431 n10__i5__i6__i2__net22 vss 73.2439e-18
c5432 n1750__chipdriverout vss 282.935e-18
c5433 n4__i5__i6__i2__net21 vss 665.891e-21
c5434 n5__i5__i7__i7__net3 vss 99.8184e-21
c5435 n1711__chipdriverout vss 415.753e-18
c5436 n8__i5__i6__net30 vss 35.19e-18
c5437 n5__i5__r2 vss 60.3588e-18
c5438 n284__vdd vss 74.1694e-18
c5439 n10__i5__i6__net30 vss 152.204e-18
c5440 n965__vddio vss 426.504e-18
c5441 n3__i5__r2 vss 70.0245e-18
c5442 n1658__chipdriverout vss 372.799e-18
c5443 n12__i5__i6__net30 vss 182.067e-18
c5444 n43__vdd vss 50.882e-18
c5445 n944__vddio vss 416.824e-18
c5446 n5__i5__i7__i7__net2 vss 63.6342e-18
c5447 n285__vdd vss 65.1223e-18
c5448 n1619__chipdriverout vss 378.017e-18
c5449 n7__i5__i6__i6__net4 vss 99.5616e-18
c5450 n1672__chipdriverout vss 410.43e-18
c5451 n14__i5__i6__net30 vss 68.5944e-18
c5452 n45__vdd vss 47.0258e-18
c5453 n7__i5__i7__i7__net2 vss 33.0184e-18
c5454 n1633__chipdriverout vss 290.702e-18
c5455 n5__i5__i6__i6__net4 vss 166.323e-18
c5456 n338__vdd vss 62.7466e-18
c5457 n923__vddio vss 412.131e-18
c5458 n17__i5__i7__net46 vss 60.9094e-18
c5459 n1579__chipdriverout vss 271.667e-18
c5460 n13__i5__i6__net31 vss 38.9829e-18
c5461 n4__i5__r1 vss 136.152e-18
c5462 n11__i5__i6__net31 vss 40.3556e-18
c5463 n1539__chipdriverout vss 273.337e-18
c5464 n14__i5__i7__net46 vss 81.0605e-18
c5465 n1591__chipdriverout vss 365.565e-18
c5466 n8__i5__i6__net31 vss 46.5248e-18
c5467 n336__vdd vss 65.1926e-18
c5468 n892__vddio vss 413.656e-18
c5469 n14__i5__i6__net31 vss 58.6961e-18
c5470 n333__vdd vss 54.1254e-18
c5471 n1551__chipdriverout vss 364.166e-18
c5472 n20__i5__i7__i7__net1 vss 62.725e-18
c5473 n884__vddio vss 410.549e-18
c5474 n21__i5__i7__net50 vss 75.4001e-18
c5475 n6__i5__i7__i7__i1__net1 vss 169.657e-18
c5476 n24__i5__i7__net50 vss 65.4079e-18
c5477 n1511__chipdriverout vss 389.918e-18
c5478 n4__i5__r0 vss 140.119e-18
c5479 n3__i5__i7__i7__i1__net1 vss 86.4558e-18
c5480 n286__vdd vss 62.9051e-18
c5481 n850__vddio vss 416.607e-18
c5482 n1499__chipdriverout vss 271.666e-18
c5483 n7__i5__r0 vss 139.572e-18
c5484 n4__i5__i7__i7__i1__net1 vss 108.807e-18
c5485 n22__i5__i7__net51 vss 58.5936e-18
c5486 n1478__chipdriverout vss 390.659e-18
c5487 n13__i5__i7__i6__net1 vss 154.729e-18
c5488 n1472__chipdriverout vss 405.693e-18
c5489 n842__vddio vss 419.2e-18
c5490 n13__i5__i7__net44 vss 21.4522e-21
c5491 n1417__chipdriverout vss 364.24e-18
c5492 n9__i5__i7__i7__net1 vss 148.573e-18
c5493 n6__i5__i7__net46 vss 67.1777e-18
c5494 n802__vddio vss 413.859e-18
c5495 n10__i5__i7__net50 vss 104.942e-21
c5496 n13__i5__i7__net47 vss 60.0149e-18
c5497 n1378__chipdriverout vss 363.692e-18
c5498 n12__i5__i7__net50 vss 19.2632e-21
c5499 n17__i5__i7__net44 vss 64.0707e-18
c5500 n7__i5__i7__net46 vss 69.4551e-18
c5501 n1405__chipdriverout vss 270.408e-18
c5502 n12__i5__i7__i7__net1 vss 135.981e-18
c5503 n6__i5__i7__i7__i0__net1 vss 172.237e-18
c5504 n1366__chipdriverout vss 271.398e-18
c5505 n777__vddio vss 403.303e-18
c5506 n3__i5__i7__i7__i0__net1 vss 89.3868e-18
c5507 n9__i5__i7__i6__net1 vss 63.4143e-18
c5508 n1339__chipdriverout vss 369.741e-18
c5509 n287__vdd vss 64.588e-18
c5510 n327__vdd vss 60.0956e-18
c5511 n4__i5__i7__i7__i0__net1 vss 109.791e-18
c5512 n11__i5__i7__i6__net1 vss 25.8405e-18
c5513 n1327__chipdriverout vss 276.977e-18
c5514 n756__vddio vss 409.999e-18
c5515 n1300__chipdriverout vss 377.3e-18
c5516 n23__i5__i7__xor3 vss 77.3574e-18
c5517 n23__i5__i7__xor0 vss 67.6152e-18
c5518 n735__vddio vss 428.009e-18
c5519 n8__i5__i7__net51 vss 149.569e-18
c5520 n4__i5__i7__net50 vss 141.327e-18
c5521 n1261__chipdriverout vss 378.506e-18
c5522 n714__vddio vss 411.323e-18
c5523 n22__i5__i7__xor2 vss 56.8957e-18
c5524 n22__i5__i7__xor1 vss 56.8306e-18
c5525 n1288__chipdriverout vss 286.822e-18
c5526 n221__vdd vss 415.063e-18
c5527 n322__vdd vss 649.187e-18
c5528 n26__i5__i7__xor3 vss 64.6191e-18
c5529 n26__i5__i7__xor0 vss 59.9734e-18
c5530 n11__i5__i7__net51 vss 139.947e-18
c5531 n7__i5__i7__net50 vss 139.114e-18
c5532 n1249__chipdriverout vss 285.848e-18
c5533 n13__i5__i7__i5__net1 vss 153.389e-18
c5534 n13__i5__i7__i4__net1 vss 155.115e-18
c5535 n1222__chipdriverout vss 389.512e-18
c5536 n693__vddio vss 400.093e-18
c5537 n8__i5__i7__net47 vss 71.8709e-18
c5538 n6__i5__i7__net44 vss 68.0974e-18
c5539 n1183__chipdriverout vss 373.625e-18
c5540 n10__i5__i7__xor3 vss 40.2256e-21
c5541 n10__i5__i7__xor0 vss 104.942e-21
c5542 n685__vddio vss 411.789e-18
c5543 n1210__chipdriverout vss 411.468e-18
c5544 n12__i5__i7__xor3 vss 12.0854e-21
c5545 n12__i5__i7__xor0 vss 19.1826e-21
c5546 n9__i5__i7__net47 vss 70.6816e-18
c5547 n7__i5__i7__net44 vss 71.2113e-18
c5548 n1171__chipdriverout vss 274.276e-18
c5549 n1132__chipdriverout vss 282.93e-18
c5550 n9__i5__i7__i5__net1 vss 26.4295e-18
c5551 n9__i5__i7__i4__net1 vss 26.3573e-18
c5552 n1119__chipdriverout vss 291.94e-18
c5553 n1144__chipdriverout vss 368.323e-18
c5554 n651__vddio vss 422.016e-18
c5555 n7__i5__i7__i5__net1 vss 64.6948e-18
c5556 n7__i5__i7__i4__net1 vss 62.5361e-18
c5557 n288__vdd vss 59.1915e-18
c5558 n321__vdd vss 62.3238e-18
c5559 n1125__chipdriverout vss 385.071e-18
c5560 n620__vddio vss 415.336e-18
c5561 n1066__chipdriverout vss 389.56e-18
c5562 n14__i5__i7__x3out vss 75.3361e-18
c5563 n14__i5__i7__x0out vss 71.3877e-18
c5564 n4__i5__i7__xor3 vss 143.661e-18
c5565 n4__i5__i7__xor0 vss 139.011e-18
c5566 n612__vddio vss 405.131e-18
c5567 n1027__chipdriverout vss 368.271e-18
c5568 n15__i5__i7__y3out vss 61.1359e-18
c5569 n17__i5__i7__y0out vss 61.1149e-18
c5570 n578__vddio vss 411.409e-18
c5571 n1054__chipdriverout vss 283.306e-18
c5572 n228__vdd vss 269.064e-18
c5573 n317__vdd vss 320.19e-18
c5574 n17__i5__i7__x3out vss 65.6669e-18
c5575 n17__i5__i7__x0out vss 66.1788e-18
c5576 n7__i5__i7__xor3 vss 135.663e-18
c5577 n7__i5__i7__xor0 vss 135.717e-18
c5578 n1015__chipdriverout vss 266.611e-18
c5579 n6__i5__i7__i9__net1 vss 170.612e-18
c5580 n6__i5__i7__i2__net1 vss 171.616e-18
c5581 n1008__chipdriverout vss 399.083e-18
c5582 n3__i5__i7__i9__net1 vss 89.304e-18
c5583 n3__i5__i7__i2__net1 vss 86.504e-18
c5584 n289__vdd vss 62.7664e-18
c5585 n316__vdd vss 61.9654e-18
c5586 n560__vddio vss 422.288e-18
c5587 n1002__chipdriverout vss 410.667e-18
c5588 n4__i5__i7__i9__net1 vss 109.149e-18
c5589 n4__i5__i7__i2__net1 vss 112.418e-18
c5590 n949__chipdriverout vss 381.091e-18
c5591 n526__vddio vss 412.276e-18
c5592 n14__i5__i7__x2out vss 76.7543e-18
c5593 n14__i5__i7__x1out vss 73.1198e-18
c5594 n910__chipdriverout vss 358.32e-18
c5595 n4__i5__i7__xor2 vss 143.248e-18
c5596 n4__i5__i7__xor1 vss 139.59e-18
c5597 n505__vddio vss 413.336e-18
c5598 n17__i5__i7__y2out vss 60.5788e-18
c5599 n17__i5__i7__y1out vss 60.7919e-18
c5600 n860__chipdriverout vss 383.603e-18
c5601 n937__chipdriverout vss 267.146e-18
c5602 n233__vdd vss 253.277e-18
c5603 n312__vdd vss 384.838e-18
c5604 n17__i5__i7__x2out vss 63.3861e-18
c5605 n17__i5__i7__x1out vss 63.4632e-18
c5606 n898__chipdriverout vss 282.778e-18
c5607 n7__i5__i7__xor2 vss 135.95e-18
c5608 n7__i5__i7__xor1 vss 135.847e-18
c5609 n6__i5__i7__i8__net1 vss 169.551e-18
c5610 n6__i5__i7__i3__net1 vss 169.705e-18
c5611 n882__chipdriverout vss 267.082e-18
c5612 n484__vddio vss 430.302e-18
c5613 n3__i5__i7__i8__net1 vss 92.1577e-18
c5614 n3__i5__i7__i3__net1 vss 90.1469e-18
c5615 n832__chipdriverout vss 390.797e-18
c5616 n290__vdd vss 65.1018e-18
c5617 n311__vdd vss 63.0393e-18
c5618 n4__i5__i7__i8__net1 vss 114.109e-18
c5619 n4__i5__i7__i3__net1 vss 111.859e-18
c5620 n820__chipdriverout vss 272.985e-18
c5621 n463__vddio vss 418.99e-18
c5622 n793__chipdriverout vss 390.21e-18
c5623 n449__vddio vss 418.614e-18
c5624 n8__i5__i7__y3out vss 74.4468e-18
c5625 n6__i5__i7__x3out vss 65.6008e-18
c5626 n743__chipdriverout vss 375.172e-18
c5627 n428__vddio vss 409.64e-18
c5628 n2__i5__i7__i1__i2__net24 vss 49.622e-18
c5629 n2__i5__i7__i0__i2__net24 vss 49.8721e-18
c5630 n291__vdd vss 64.4122e-18
c5631 n308__vdd vss 64.6307e-18
c5632 n704__chipdriverout vss 404.335e-18
c5633 n5__i5__i7__i1__i2__net22 vss 45.6011e-18
c5634 n5__i5__i7__i0__i2__net22 vss 44.2638e-18
c5635 n403__vddio vss 413.131e-18
c5636 n665__chipdriverout vss 371.547e-18
c5637 n2__i5__i7__i1__i2__net21 vss 50.2759e-18
c5638 n2__i5__i7__i0__i2__net21 vss 47.536e-18
c5639 n382__vddio vss 404.44e-18
c5640 n292__vdd vss 63.9301e-18
c5641 n307__vdd vss 64.0141e-18
c5642 n6__i5__i7__y3out vss 111.695e-18
c5643 n4__i5__i7__x3out vss 112.565e-18
c5644 n781__chipdriverout vss 267.956e-18
c5645 n237__vdd vss 1.25154e-15
c5646 n256__vdd vss 1.62284e-15
c5647 n10__i5__i7__y3out vss 54.2415e-18
c5648 n8__i5__i7__x3out vss 53.7228e-18
c5649 n757__chipdriverout vss 384.632e-18
c5650 n2__i5__i7__i1__i2__net25 vss 32.8185e-18
c5651 n2__i5__i7__i0__i2__net25 vss 33.6735e-18
c5652 n718__chipdriverout vss 277.311e-18
c5653 n7__i5__i7__i1__i2__net22 vss 31.2322e-18
c5654 n7__i5__i7__i0__i2__net22 vss 31.0606e-18
c5655 n679__chipdriverout vss 281.158e-18
c5656 n2__i5__i7__i1__i2__net23 vss 31.7305e-18
c5657 n2__i5__i7__i0__i2__net23 vss 32.1481e-18
c5658 n640__chipdriverout vss 271.673e-18
c5659 n4__i5__i7__y2out vss 111.282e-18
c5660 n4__i5__i7__x2out vss 112.372e-18
c5661 n601__chipdriverout vss 271.041e-18
c5662 n8__i5__i7__y2out vss 54.8185e-18
c5663 n8__i5__i7__x2out vss 54.3417e-18
c5664 n2__i5__i7__i1__i1__net25 vss 33.5542e-18
c5665 n2__i5__i7__i0__i1__net25 vss 34.2216e-18
c5666 n580__chipdriverout vss 271.223e-18
c5667 n7__i5__i7__i1__i1__net22 vss 31.6606e-18
c5668 n7__i5__i7__i0__i1__net22 vss 31.5987e-18
c5669 n541__chipdriverout vss 401.81e-18
c5670 n2__i5__i7__i1__i1__net23 vss 31.4188e-18
c5671 n2__i5__i7__i0__i1__net23 vss 31.3845e-18
c5672 n484__chipdriverout vss 271.384e-18
c5673 n626__chipdriverout vss 370.345e-18
c5674 n361__vddio vss 414.157e-18
c5675 n587__chipdriverout vss 392.409e-18
c5676 n6__i5__i7__y2out vss 72.5365e-18
c5677 n6__i5__i7__x2out vss 68.289e-18
c5678 n327__vddio vss 418.119e-18
c5679 n2__i5__i7__i1__i1__net24 vss 50.1255e-18
c5680 n2__i5__i7__i0__i1__net24 vss 51.1792e-18
c5681 n573__chipdriverout vss 394.149e-18
c5682 n293__vdd vss 64.9049e-18
c5683 n306__vdd vss 66.6267e-18
c5684 n319__vddio vss 408.594e-18
c5685 n5__i5__i7__i1__i1__net22 vss 47.2162e-18
c5686 n5__i5__i7__i0__i1__net22 vss 45.2378e-18
c5687 n534__chipdriverout vss 371.039e-18
c5688 n285__vddio vss 403.935e-18
c5689 n2__i5__i7__i1__i1__net21 vss 50.5256e-18
c5690 n2__i5__i7__i0__i1__net21 vss 47.4724e-18
c5691 n294__vdd vss 63.862e-18
c5692 n305__vdd vss 65.5376e-18
c5693 n470__chipdriverout vss 365.361e-18
c5694 n430__chipdriverout vss 292.7e-18
c5695 n5__i5__i7__y1out vss 54.5703e-18
c5696 n5__i5__i7__x1out vss 54.6317e-18
c5697 n391__chipdriverout vss 282.099e-18
c5698 n2__i5__i7__i1__i0__net25 vss 33.4507e-18
c5699 n2__i5__i7__i0__i0__net25 vss 33.8561e-18
c5700 n7__i5__i7__i1__i0__net22 vss 31.6796e-18
c5701 n7__i5__i7__i0__i0__net22 vss 32.3434e-18
c5702 n352__chipdriverout vss 282.265e-18
c5703 n2__i5__i7__i1__i0__net23 vss 31.7062e-18
c5704 n2__i5__i7__i0__i0__net23 vss 31.5706e-18
c5705 n313__chipdriverout vss 283.169e-18
c5706 n254__vddio vss 398.517e-18
c5707 n442__chipdriverout vss 412.5e-18
c5708 n3__i5__i7__y1out vss 72.0375e-18
c5709 n3__i5__i7__x1out vss 69.3392e-18
c5710 n246__vddio vss 426.746e-18
c5711 n403__chipdriverout vss 390.797e-18
c5712 n2__i5__i7__i1__i0__net24 vss 49.6005e-18
c5713 n2__i5__i7__i0__i0__net24 vss 52.1328e-18
c5714 n295__vdd vss 63.4183e-18
c5715 n304__vdd vss 67.5215e-18
c5716 n212__vddio vss 411.15e-18
c5717 n5__i5__i7__i1__i0__net22 vss 45.0452e-18
c5718 n5__i5__i7__i0__i0__net22 vss 46.6824e-18
c5719 n364__chipdriverout vss 366.471e-18
c5720 n181__vddio vss 404.42e-18
c5721 n2__i5__i7__i1__i0__net21 vss 50.6783e-18
c5722 n2__i5__i7__i0__i0__net21 vss 48.6076e-18
c5723 n325__chipdriverout vss 367.84e-18
c5724 n296__vdd vss 63.1857e-18
c5725 n303__vdd vss 64.8616e-18
c5726 n274__chipdriverout vss 410.868e-18
c5727 n5__i5__i7__y0out vss 52.5969e-18
c5728 n5__i5__i7__x0out vss 54.9604e-18
c5729 n235__chipdriverout vss 282.2e-18
c5730 n2__i5__i7__i1__i3__net25 vss 33.7895e-18
c5731 n2__i5__i7__i0__i3__net25 vss 33.632e-18
c5732 n196__chipdriverout vss 273.917e-18
c5733 n7__i5__i7__i1__i3__net22 vss 31.3299e-18
c5734 n7__i5__i7__i0__i3__net22 vss 32.5904e-18
c5735 n157__chipdriverout vss 272.749e-18
c5736 n2__i5__i7__i1__i3__net23 vss 35.6544e-18
c5737 n2__i5__i7__i0__i3__net23 vss 35.7369e-18
c5738 n160__vddio vss 408.967e-18
c5739 n286__chipdriverout vss 392.082e-18
c5740 n139__vddio vss 414.802e-18
c5741 n3__i5__i7__y0out vss 79.5452e-18
c5742 n3__i5__i7__x0out vss 75.2674e-18
c5743 n247__chipdriverout vss 390.426e-18
c5744 n2__i5__i7__i1__i3__net24 vss 50.5838e-18
c5745 n2__i5__i7__i0__i3__net24 vss 51.2339e-18
c5746 n118__vddio vss 409.945e-18
c5747 n297__vdd vss 66.7438e-18
c5748 n302__vdd vss 66.5964e-18
c5749 n208__chipdriverout vss 363.291e-18
c5750 n5__i5__i7__i1__i3__net22 vss 45.4368e-18
c5751 n5__i5__i7__i0__i3__net22 vss 45.4145e-18
c5752 n97__vddio vss 409.389e-18
c5753 n169__chipdriverout vss 368.11e-18
c5754 n2__i5__i7__i1__i3__net21 vss 52.7063e-18
c5755 n2__i5__i7__i0__i3__net21 vss 50.8328e-18
c5756 n298__vdd vss 68.4483e-18
c5757 n301__vdd vss 69.6154e-18
c5758 n70__vddio vss 429.424e-18
c5759 n8__i5__i7__i1__net1 vss 46.7947e-18
c5760 n133__chipdriverout vss 272.195e-18
c5761 n8__i5__i7__i0__net1 vss 44.8468e-18
c5762 n9__i5__i7__i1__net1 vss 62.9659e-18
c5763 n119__chipdriverout vss 390.498e-18
c5764 n9__i5__i7__i0__net1 vss 62.6311e-18
c5765 n299__vdd vss 56.4723e-18
c5766 n300__vdd vss 64.7393e-18
c5767 n45__vddio vss 418.059e-18
c5768 n80__chipdriverout vss 390.498e-18
c5769 n24__vddio vss 417.929e-18
c5770 n41__chipdriverout vss 392.701e-18
c5771 n3__vddio vss 416.681e-18
c5772 n3__chipdriverout vss 274.463e-18
c5773 n94__chipdriverout vss 272.067e-18
c5774 n55__chipdriverout vss 409.607e-18
c5775 n16__chipdriverout vss 195.585e-18
c5776 n2__x0 vss 15.7705e-18
c5777 n2__y0 vss 15.9756e-18
c5778 n2__i5__i7__i0__i3__net22 vss 15.0704e-18
c5779 n2__i5__i7__i1__i3__net22 vss 15.8349e-18
c5780 n17__chipdriverout vss 64.1291e-18
c5781 n2__x1 vss 16.3188e-18
c5782 n2__y1 vss 16.4992e-18
c5783 n56__chipdriverout vss 85.7296e-18
c5784 n95__chipdriverout vss 84.6606e-18
c5785 n2__i5__i7__i0__i0__net22 vss 15.0805e-18
c5786 n2__i5__i7__i1__i0__net22 vss 15.8798e-18
c5787 n134__chipdriverout vss 84.5238e-18
c5788 n158__chipdriverout vss 84.5127e-18
c5789 n197__chipdriverout vss 84.6503e-18
c5790 n6__i5__i7__i0__i3__net22 vss 33.8221e-18
c5791 n6__i5__i7__i1__i3__net22 vss 33.9777e-18
c5792 n2__x2 vss 16.7419e-18
c5793 n2__y2 vss 15.6285e-18
c5794 n236__chipdriverout vss 83.0614e-18
c5795 n2__i5__i7__i0__i1__net22 vss 15.6538e-18
c5796 n2__i5__i7__i1__i1__net22 vss 15.7093e-18
c5797 n275__chipdriverout vss 83.5394e-18
c5798 n314__chipdriverout vss 83.0283e-18
c5799 n353__chipdriverout vss 83.1678e-18
c5800 n2__x3 vss 15.6354e-18
c5801 n6__i5__i7__i0__i0__net22 vss 35.2484e-18
c5802 n6__i5__i7__i1__i0__net22 vss 35.9079e-18
c5803 n2__y3 vss 16.9413e-18
c5804 n392__chipdriverout vss 83.0614e-18
c5805 n431__chipdriverout vss 88.2826e-18
c5806 n2__i5__i7__i0__i2__net22 vss 14.646e-18
c5807 n2__i5__i7__i1__i2__net22 vss 15.7332e-18
c5808 n485__chipdriverout vss 84.4619e-18
c5809 n8__x2 vss 29.9284e-18
c5810 n9__x2 vss 22.4789e-18
c5811 n542__chipdriverout vss 84.6509e-18
c5812 n6__i5__i7__i0__i1__net22 vss 36.2763e-18
c5813 n6__i5__i7__i1__i1__net22 vss 36.8324e-18
c5814 n581__chipdriverout vss 84.4272e-18
c5815 n602__chipdriverout vss 84.9206e-18
c5816 n641__chipdriverout vss 83.7545e-18
c5817 n7__x3 vss 30.6747e-18
c5818 n8__x3 vss 25.5935e-18
c5819 n680__chipdriverout vss 84.4385e-18
c5820 n719__chipdriverout vss 84.4109e-18
c5821 n6__i5__i7__i0__i2__net22 vss 35.9665e-18
c5822 n6__i5__i7__i1__i2__net22 vss 37.0267e-18
c5823 n758__chipdriverout vss 76.4277e-18
c5824 n782__chipdriverout vss 86.2358e-18
c5825 n821__chipdriverout vss 85.2113e-18
c5826 n883__chipdriverout vss 86.3663e-18
c5827 n899__chipdriverout vss 85.834e-18
c5828 n15__i5__i7__x2out vss 81.8792e-18
c5829 n15__i5__i7__x1out vss 77.2446e-18
c5830 n938__chipdriverout vss 86.4612e-18
c5831 n1003__chipdriverout vss 85.8257e-18
c5832 n1016__chipdriverout vss 89.4447e-18
c5833 n15__i5__i7__x3out vss 86.5244e-18
c5834 n15__i5__i7__x0out vss 85.8187e-18
c5835 n1055__chipdriverout vss 83.3601e-18
c5836 n1120__chipdriverout vss 83.5506e-18
c5837 n1133__chipdriverout vss 83.3943e-18
c5838 n8__i5__i7__i5__net1 vss 87.6334e-18
c5839 n8__i5__i7__i4__net1 vss 88.5787e-18
c5840 n1172__chipdriverout vss 83.8944e-18
c5841 n20__i5__i7__xor2 vss 309.603e-18
c5842 n20__i5__i7__xor1 vss 264.716e-18
c5843 n14__i5__i7__xor3 vss 41.1071e-18
c5844 n14__i5__i7__xor0 vss 41.2863e-18
c5845 n16__i5__i7__xor0 vss 42.1017e-18
c5846 n1211__chipdriverout vss 83.4042e-18
c5847 n19__i5__i7__xor3 vss 206.764e-18
c5848 n21__i5__i7__xor3 vss 126.193e-18
c5849 n19__i5__i7__xor0 vss 207.158e-18
c5850 n21__i5__i7__xor0 vss 123.648e-18
c5851 n1250__chipdriverout vss 83.501e-18
c5852 n21__i5__i7__xor2 vss 114.449e-18
c5853 n21__i5__i7__xor1 vss 111.098e-18
c5854 n24__i5__i7__xor3 vss 95.4856e-18
c5855 n24__i5__i7__xor0 vss 95.6951e-18
c5856 n2__i5__clk_buf vss 12.4461e-18
c5857 n7__i5__clk_buf vss 11.4649e-18
c5858 n1289__chipdriverout vss 83.3601e-18
c5859 n1328__chipdriverout vss 83.7808e-18
c5860 n1367__chipdriverout vss 84.2576e-18
c5861 n10__i5__i7__i6__net1 vss 88.7329e-18
c5862 n1406__chipdriverout vss 83.4832e-18
c5863 n15__i5__i7__net44 vss 90.5036e-18
c5864 n14__i5__i7__net50 vss 41.2577e-18
c5865 n16__i5__i7__net50 vss 42.0934e-18
c5866 n20__i5__i7__net51 vss 197.634e-18
c5867 n2__i5__i6__net30 vss 6.44813e-18
c5868 n4__i5__i6__net30 vss 6.82167e-18
c5869 n19__i5__i7__net50 vss 208.304e-18
c5870 n2__i5__i6__net31 vss 15.7873e-18
c5871 n1473__chipdriverout vss 84.6143e-18
c5872 n1500__chipdriverout vss 84.14e-18
c5873 n21__i5__i7__net51 vss 116.571e-18
c5874 n2__i5__i6__i2__net22 vss 6.54217e-18
c5875 n4__i5__i6__i2__net22 vss 7.46863e-18
c5876 n22__i5__i7__net50 vss 100.23e-18
c5877 n1540__chipdriverout vss 84.3106e-18
c5878 n37__reset vss 16.7601e-18
c5879 n15__i5__i7__net46 vss 84.6268e-18
c5880 n1580__chipdriverout vss 84.1234e-18
c5881 n9__i5__i6__net31 vss 36.2675e-18
c5882 n10__i5__i6__net31 vss 67.3958e-18
c5883 n24__i5__i7__i7__net1 vss 117.828e-18
c5884 n25__i5__i7__i7__net1 vss 73.9648e-18
c5885 n1634__chipdriverout vss 87.8986e-18
c5886 n1673__chipdriverout vss 83.4081e-18
c5887 n75__vdd vss 49.3729e-18
c5888 n86__vdd vss 18.6542e-18
c5889 n88__vdd vss 12.2034e-18
c5890 n94__vdd vss 17.0857e-18
c5891 n108__vdd vss 11.0491e-18
c5892 n114__vdd vss 11.0001e-18
c5893 n116__vdd vss 7.28671e-18
c5894 n127__vdd vss 20.146e-18
c5895 n133__vdd vss 21.253e-18
c5896 n135__vdd vss 22.8321e-18
c5897 n141__vdd vss 22.9883e-18
c5898 n1712__chipdriverout vss 83.6247e-18
c5899 n6__i5__i7__i7__net2 vss 81.6851e-18
c5900 n8__i5__i7__i7__net2 vss 125.518e-18
c5901 n19__i5__clk_buf vss 12.9938e-18
c5902 n24__i5__clk_buf vss 11.8157e-18
c5903 n6__i5__i7__i7__net3 vss 142.824e-18
c5904 n20__i5__i7__net46 vss 214.566e-18
c5905 n21__i5__i7__net46 vss 305.446e-18
c5906 n2__i5__i6__net33 vss 6.43994e-18
c5907 n4__i5__i6__net33 vss 6.81779e-18
c5908 n1751__chipdriverout vss 83.4035e-18
c5909 n19__i5__i6__net31 vss 15.7218e-18
c5910 n2__i5__i8__net1 vss 8.4132e-18
c5911 n4__i5__i8__net1 vss 9.52861e-18
c5912 n9__i5__i6__i2__net21 vss 44.8513e-18
c5913 n1790__chipdriverout vss 83.8848e-18
c5914 n2__i5__i8__net4 vss 15.3667e-18
c5915 n9__i5__i6__i2__net22 vss 78.7967e-18
c5916 n2__i5__i6__i4__net22 vss 6.28218e-18
c5917 n4__i5__i6__i4__net22 vss 7.4617e-18
c5918 n25__i5__i6__net31 vss 107.685e-18
c5919 n9__i5__i6__i2__net23 vss 32.9756e-18
c5920 n1824__chipdriverout vss 83.4017e-18
c5921 n2__i5__i8__i9__net22 vss 8.78136e-18
c5922 n4__i5__i8__i9__net22 vss 7.59833e-18
c5923 n1868__chipdriverout vss 83.5104e-18
c5924 n44__reset vss 16.7651e-18
c5925 n3__i5__i6__net32 vss 41.8782e-18
c5926 n4__i5__i6__net32 vss 56.8227e-18
c5927 n153__vdd vss 25.7644e-18
c5928 n19__i5__i9__net21 vss 86.9936e-18
c5929 n48__reset vss 12.9813e-18
c5930 n1907__chipdriverout vss 84.2165e-18
c5931 n2__i5__i8__net2 vss 13.874e-18
c5932 n7__i5__i8__net2 vss 12.5107e-18
c5933 n45__i5__clk_buf vss 77.3212e-18
c5934 n46__i5__clk_buf vss 82.7262e-18
c5935 n2__i5__i6__net35 vss 5.8469e-18
c5936 n4__i5__i6__net35 vss 6.8122e-18
c5937 n2__i5__i8__net5 vss 8.56822e-18
c5938 n4__i5__i8__net5 vss 7.14611e-18
c5939 n9__i5__i8__net4 vss 35.7752e-18
c5940 n10__i5__i8__net4 vss 74.4755e-18
c5941 n9__i5__i6__i4__net21 vss 46.3759e-18
c5942 n33__i5__i6__net31 vss 15.7746e-18
c5943 n12__i5__i8__net1 vss 16.6395e-18
c5944 n793__i1__i14__net1 vss 84.7605e-18
c5945 n9__i5__i6__i4__net22 vss 78.9797e-18
c5946 n9__i5__i8__i9__net21 vss 43.3955e-18
c5947 n2__i5__i6__i5__net22 vss 5.48189e-18
c5948 n4__i5__i6__i5__net22 vss 7.95326e-18
c5949 n2__i5__i8__i10__net22 vss 7.3387e-18
c5950 n4__i5__i8__i10__net22 vss 7.67926e-18
c5951 n37__i5__i6__net31 vss 109.209e-18
c5952 n9__i5__i6__i4__net23 vss 34.0027e-18
c5953 n832__i1__i14__net1 vss 83.4819e-18
c5954 n9__i5__i8__i9__net22 vss 79.5507e-18
c5955 n17__i5__i8__net4 vss 220.02e-18
c5956 n7__i5__i8__i9__net23 vss 34.4954e-18
c5957 n871__i1__i14__net1 vss 84.6239e-18
c5958 n3__i5__i6__net34 vss 42.5327e-18
c5959 n4__i5__i6__net34 vss 57.3428e-18
c5960 n57__reset vss 15.9849e-18
c5961 n61__reset vss 10.9853e-18
c5962 n66__reset vss 1.53476e-15
c5963 n910__i1__i14__net1 vss 84.1325e-18
c5964 n77__i5__clk4 vss 11.4606e-18
c5965 n82__i5__clk4 vss 13.0065e-18
c5966 n20__i5__i8__net2 vss 19.5056e-18
c5967 n21__i5__i8__net2 vss 9.20574e-18
c5968 n22__i5__i8__net2 vss 41.8228e-18
c5969 n23__i5__i8__net2 vss 36.0848e-18
c5970 n24__i5__i8__net2 vss 56.1731e-18
c5971 n949__i1__i14__net1 vss 84.3483e-18
c5972 n86__i5__clk4 vss 21.7316e-18
c5973 n20__i5__i8__net1 vss 55.5651e-18
c5974 n988__i1__i14__net1 vss 84.11e-18
c5975 n2__piso_out vss 23.3456e-18
c5976 n3__piso_out vss 15.9903e-18
c5977 n4__piso_out vss 14.1214e-18
c5978 n5__piso_out vss 18.4668e-18
c5979 n1042__i1__i14__net1 vss 87.9089e-18
c5980 n7__i5__i6__i5__net21 vss 45.3991e-18
c5981 n7__i5__i8__i10__net21 vss 59.5042e-18
c5982 n1099__i1__i14__net1 vss 83.4891e-18
c5983 n9__i5__i6__i5__net22 vss 80.1915e-18
c5984 n9__i5__i8__i10__net22 vss 80.9835e-18
c5985 n45__i5__i6__net31 vss 110.42e-18
c5986 n1105__i1__i14__net1 vss 83.5245e-18
c5987 n7__i5__i6__i5__net23 vss 33.0637e-18
c5988 n69__i5__clk_buf vss 285.772e-18
c5989 n70__i5__clk_buf vss 228.162e-18
c5990 n71__i5__clk_buf vss 258.823e-18
c5991 n9__i5__i8__i10__net23 vss 34.758e-18
c5992 n46__i5__i6__net31 vss 408.169e-18
c5993 n47__i5__i6__net31 vss 396.986e-18
c5994 n1144__i1__i14__net1 vss 83.4035e-18
c5995 n5__bufin vss 34.8925e-18
c5996 n6__bufin vss 42.7772e-18
c5997 n7__bufin vss 58.4712e-18
c5998 n1198__i1__i14__net1 vss 83.8944e-18
c5999 n89__i5__clk4 vss 23.7518e-18
c6000 n90__i5__clk4 vss 26.8183e-18
c6001 n91__i5__clk4 vss 47.1204e-18
c6002 n92__i5__clk4 vss 64.0844e-18
c6003 n8__i4__net1 vss 57.3779e-18
c6004 n14__i5__i8__net5 vss 43.7315e-18
c6005 n15__i5__i8__net5 vss 62.4008e-18
c6006 n1237__i1__i14__net1 vss 83.395e-18
c6007 n15__piso_out vss 61.4739e-18
c6008 n1261__i1__i14__net1 vss 83.5097e-18
c6009 n42__shift vss 1.14874e-15
c6010 n43__shift vss 525.696e-18
c6011 n5__piso_outinv vss 63.1437e-18
c6012 n5__i5__i8__i8__net1 vss 58.3412e-18
c6013 n1326__i1__i14__net1 vss 84.2254e-18
c6014 n185__vdd vss 164.21e-18
c6015 n191__vdd vss 374.159e-18
c6016 n196__vdd vss 292.343e-18
c6017 n199__vdd vss 48.9077e-18
c6018 n200__vdd vss 36.4341e-18
c6019 n202__vdd vss 32.5083e-18
c6020 n205__vdd vss 140.031e-18
c6021 n206__vdd vss 32.1152e-18
c6022 n208__vdd vss 61.6397e-18
c6023 n209__vdd vss 61.4346e-18
c6024 n211__vdd vss 58.4692e-18
c6025 n220__vdd vss 111.569e-18
c6026 n226__vdd vss 63.3169e-18
c6027 n231__vdd vss 68.4624e-18
c6028 n236__vdd vss 76.3903e-18
c6029 n241__vdd vss 65.8424e-18
c6030 n245__vdd vss 58.5543e-18
c6031 n254__vdd vss 194.535e-18
c6032 n255__vdd vss 157.389e-18
c6033 n258__vdd vss 76.1607e-18
c6034 n261__vdd vss 80.9994e-18
c6035 n264__vdd vss 76.5003e-18
c6036 n267__vdd vss 77.2812e-18
c6037 n310__vdd vss 39.1478e-18
c6038 n315__vdd vss 129.404e-18
c6039 n320__vdd vss 55.1553e-18
c6040 n326__vdd vss 69.7746e-18
c6041 n332__vdd vss 63.0291e-18
c6042 n337__vdd vss 35.51e-18
c6043 n340__vdd vss 148.609e-18
c6044 n343__vdd vss 109.001e-18
c6045 n346__vdd vss 56.3177e-18
c6046 n349__vdd vss 154.807e-18
c6047 n352__vdd vss 107.875e-18
c6048 n355__vdd vss 55.2844e-18
c6049 n358__vdd vss 153.987e-18
c6050 n361__vdd vss 114.811e-18
c6051 n364__vdd vss 34.1101e-18
c6052 n369__vdd vss 28.186e-18
c6053 n371__vdd vss 32.3065e-18
c6054 n376__vdd vss 27.4822e-18
c6055 n380__vdd vss 57.56e-18
c6056 n1531__vddio vss 3.23852e-18
c6057 n1532__vddio vss 1.7382e-18
c6058 n1535__vddio vss 3.66701e-18
c6059 n1536__vddio vss 3.69039e-18
c6060 n1537__vddio vss 1.81341e-18
c6061 n1540__vddio vss 3.80722e-18
c6062 n1541__vddio vss 3.66012e-18
c6063 n1542__vddio vss 1.64206e-18
c6064 n1545__vddio vss 3.23988e-18
c6065 n1546__vddio vss 2.01145e-18
c6066 n1549__vddio vss 1.68203e-18
c6067 n1550__vddio vss 3.68353e-18
c6068 n1553__vddio vss 3.44775e-18
c6069 n1554__vddio vss 3.54329e-18
c6070 n1557__vddio vss 3.52422e-18
c6071 n1558__vddio vss 3.6835e-18
c6072 n1561__vddio vss 3.46973e-18
c6073 n1562__vddio vss 3.12304e-18
c6074 n1565__vddio vss 3.67336e-18
c6075 n1566__vddio vss 3.57516e-18
c6076 n1569__vddio vss 3.23162e-18
c6077 n1570__vddio vss 3.51145e-18
c6078 n1573__vddio vss 3.23607e-18
c6079 n1574__vddio vss 3.73205e-18
c6080 n1577__vddio vss 3.27175e-18
c6081 n1578__vddio vss 4.06827e-18
c6082 n1581__vddio vss 3.29672e-18
c6083 n1582__vddio vss 3.49955e-18
c6084 n1585__vddio vss 3.27175e-18
c6085 n1586__vddio vss 3.57145e-18
c6086 n1589__vddio vss 3.57516e-18
c6087 n1590__vddio vss 3.52979e-18
c6088 n1593__vddio vss 3.70064e-18
c6089 n1594__vddio vss 3.55274e-18
c6090 n389__vdd vss 47.933e-18
c6091 n398__vdd vss 39.6463e-18
c6092 n400__vdd vss 33.9904e-18
c6093 n20__piso_out vss 5.06569e-18
c6094 n5__i1__net3 vss 43.1285e-18
c6095 n409__vdd vss 11.3604e-18
c6096 n414__vdd vss 80.7736e-18
c6097 n418__vdd vss 53.4152e-18
c6098 n13__i1__net3 vss 64.5786e-18
c6099 n20__i1__net3 vss 71.9271e-18
c6100 n25__i1__net3 vss 65.5449e-18
c6101 n59__i1__i12__net1 vss 60.5638e-18
c6102 n60__i1__i12__net1 vss 30.9329e-18
c6103 n63__i1__i12__net1 vss 77.3226e-18
c6104 n1734__vddio vss 127.774e-18
c6105 n6__i1__i11__outinv vss 115.583e-18
c6106 n1769__vddio vss 12.9106e-18
c6107 n1773__vddio vss 18.0662e-18
c6108 n1777__vddio vss 25.6386e-18
c6109 n28__i1__net4 vss 115.709e-18
c6110 n1839__vddio vss 39.7178e-18
c6111 n79__i1__net3 vss 1.13765e-15
c6112 n215__i1__i13__net1 vss 109.407e-18
c6113 n216__i1__i13__net1 vss 22.5882e-18
c6114 n217__i1__i13__net1 vss 21.5542e-18
c6115 n218__i1__i13__net1 vss 20.8577e-18
c6116 n219__i1__i13__net1 vss 43.5462e-18
c6117 n220__i1__i13__net1 vss 18.4256e-18
c6118 n221__i1__i13__net1 vss 20.244e-18
c6119 n222__i1__i13__net1 vss 38.0354e-18
c6120 n223__i1__i13__net1 vss 37.943e-18
c6121 n224__i1__i13__net1 vss 38.1818e-18
c6122 n225__i1__i13__net1 vss 45.25e-18
c6123 n226__i1__i13__net1 vss 28.4236e-18
c6124 n84__i1__net3 vss 32.0047e-18
c6125 n1942__vddio vss 1.30738e-21
c6126 n1954__vddio vss 14.8935e-18
c6127 n1956__vddio vss 14.3053e-18
c6128 n1958__vddio vss 18.0536e-18
c6129 n1960__vddio vss 16.7897e-18
c6130 n1968__vddio vss 29.2095e-18
c6131 n1974__vddio vss 16.2906e-18
c6132 n1976__vddio vss 29.2358e-18
c6133 n1978__vddio vss 14.9247e-18
c6134 n475__vdd vss 42.7595e-18
c6135 n479__vdd vss 66.2708e-18
c6136 n2043__vddio vss 8.98394e-18
c6137 n2045__vddio vss 35.6895e-18
c6138 n2107__vddio vss 123.47e-21
c6139 n2157__vddio vss 47.8266e-18
c6140 n2156__vddio vss 3.35389e-18
rc1 chipdriverout n1577__chipdriverout 7.362e-3
rc2 n2026__vss n2039__vss 84.53e-3
rc3 n2039__vss n2015__vss 104.9e-3
rc4 n2028__vss n2039__vss 4.667e-3
rc6 n2040__vss n2042__vss 4.107e-3
rc9 n2042__vss vss 1.996e-3
rc10 vss n2045__vss 3.518e-3
rc12 n2045__vss n2019__vss 2.847e-3
rc13 n2019__vss n2047__vss 5.111e-3
rc15 n2045__vss n2049__vss 83.42e-3
rc16 n2049__vss n2050__vss 64.84e-3
rc17 n2050__vss n2051__vss 72.13e-3
rc18 n2051__vss n2052__vss 59.54e-3
rc19 n2052__vss n2053__vss 64.84e-3
rc20 n2053__vss n2054__vss 72.13e-3
rc21 n2054__vss n2055__vss 68.53e-3
rc22 n2055__vss n2056__vss 64.84e-3
rc23 n2056__vss n2057__vss 72.13e-3
rc24 n2057__vss n2058__vss 59.54e-3
rc25 n2058__vss n2059__vss 64.84e-3
rc26 n2059__vss n2060__vss 72.13e-3
rc27 n2060__vss vss 37.85e-3
rc28 vss n2061__vss 13.18e-3
rc29 vss n2062__vss 3.632e-3
rc30 n2062__vss n2063__vss 4.908e-3
rc31 n2063__vss n2064__vss 70.82e-3
rc32 n2062__vss n2065__vss 32.23e-3
rc33 n2064__vss n2066__vss 73.43e-3
rc34 n2065__vss n2067__vss 72.69e-3
rc35 n2066__vss n2068__vss 66.14e-3
rc36 n2067__vss n2069__vss 65.41e-3
rc37 n2068__vss n2070__vss 60.84e-3
rc38 n2069__vss n2071__vss 60.11e-3
rc39 n2070__vss n2072__vss 73.43e-3
rc40 n2071__vss n2073__vss 72.69e-3
rc41 n2072__vss n2074__vss 66.14e-3
rc42 n2073__vss n2075__vss 65.41e-3
rc43 n2074__vss n2076__vss 69.83e-3
rc44 n2075__vss n2077__vss 69.1e-3
rc45 n2076__vss n2078__vss 73.43e-3
rc46 n2077__vss n2079__vss 72.69e-3
rc47 n2078__vss n2080__vss 66.14e-3
rc48 n2079__vss n2081__vss 65.41e-3
rc49 n2080__vss n2082__vss 60.84e-3
rc50 n2081__vss n2083__vss 60.11e-3
rc51 n2082__vss n2084__vss 73.43e-3
rc52 n2083__vss n2085__vss 72.69e-3
rc53 n2084__vss n2086__vss 66.14e-3
rc54 n2085__vss n2087__vss 65.41e-3
rc55 n2086__vss n2088__vss 81.65e-3
rc56 n2087__vss n2089__vss 81.19e-3
rc57 n2088__vss n2040__vss 4.355e-3
rc58 n2089__vss n2042__vss 2.668e-3
rc59 n2020__vss n2040__vss 7.778e-3
rc60 n2037__vss n2040__vss 7.778e-3
rc61 n2016__vss n2042__vss 4.667e-3
rc62 n2001__vss n2042__vss 7.778e-3
rc63 n2035__vss n2042__vss 7.778e-3
rc64 n2023__vss n2045__vss 7.778e-3
rc65 n2033__vss n2045__vss 7.778e-3
rc66 n2009__vss n2047__vss 7.778e-3
rc67 n2031__vss n2047__vss 7.778e-3
rc68 n1327__vss n2049__vss 7.778e-3
rc69 n1321__vss n2050__vss 7.778e-3
rc70 n1337__vss n2051__vss 7.778e-3
rc71 n1346__vss n2052__vss 7.778e-3
rc72 n1355__vss n2053__vss 7.778e-3
rc73 n551__vss n2054__vss 7.778e-3
rc74 n1367__vss n2055__vss 7.778e-3
rc75 n1376__vss n2056__vss 7.778e-3
rc76 n1385__vss n2057__vss 7.778e-3
rc77 n1394__vss n2058__vss 7.778e-3
rc78 n1403__vss n2059__vss 7.778e-3
rc79 n1412__vss n2060__vss 7.778e-3
rc80 n1421__vss n2061__vss 7.778e-3
rc81 n1419__vss n2062__vss 7.778e-3
rc82 n1417__vss n2063__vss 7.778e-3
rc83 n1408__vss n2064__vss 7.778e-3
rc84 n1410__vss n2065__vss 7.778e-3
rc85 n1399__vss n2066__vss 7.778e-3
rc86 n1401__vss n2067__vss 7.778e-3
rc87 n1390__vss n2068__vss 7.778e-3
rc88 n1392__vss n2069__vss 7.778e-3
rc89 n1381__vss n2070__vss 7.778e-3
rc90 n1383__vss n2071__vss 7.778e-3
rc91 n1372__vss n2072__vss 7.778e-3
rc92 n1374__vss n2073__vss 7.778e-3
rc93 n1363__vss n2074__vss 7.778e-3
rc94 n1365__vss n2075__vss 7.778e-3
rc95 n547__vss n2076__vss 7.778e-3
rc96 n549__vss n2077__vss 7.778e-3
rc97 n1351__vss n2078__vss 7.778e-3
rc98 n1353__vss n2079__vss 7.778e-3
rc99 n1342__vss n2080__vss 7.778e-3
rc100 n1344__vss n2081__vss 7.778e-3
rc101 n1333__vss n2082__vss 7.778e-3
rc102 n1335__vss n2083__vss 7.778e-3
rc103 n1317__vss n2084__vss 7.778e-3
rc104 n1319__vss n2085__vss 7.778e-3
rc105 n1323__vss n2086__vss 7.778e-3
rc106 n1325__vss n2087__vss 7.778e-3
rc107 n486__vdd n487__vdd 65.52e-3
rc108 n487__vdd n488__vdd 72.8e-3
rc109 n488__vdd n489__vdd 60.21e-3
rc110 n489__vdd n490__vdd 65.52e-3
rc111 n490__vdd n491__vdd 72.8e-3
rc112 n491__vdd n492__vdd 69.21e-3
rc113 n492__vdd n493__vdd 65.52e-3
rc114 n493__vdd n494__vdd 72.8e-3
rc115 n494__vdd n495__vdd 60.21e-3
rc116 n495__vdd n496__vdd 65.52e-3
rc117 n496__vdd n497__vdd 72.8e-3
rc118 n497__vdd n498__vdd 57.71e-3
rc119 n498__vdd vdd 8.448e-3
rc120 vdd n6__vdd 5.726e-3
rc121 n6__vdd n499__vdd 68.48e-3
rc122 n499__vdd n500__vdd 72.23e-3
rc123 n500__vdd n501__vdd 64.94e-3
rc124 n501__vdd n502__vdd 59.64e-3
rc125 n502__vdd n503__vdd 72.23e-3
rc126 n503__vdd n504__vdd 64.94e-3
rc127 n504__vdd n505__vdd 68.63e-3
rc128 n505__vdd n506__vdd 72.23e-3
rc129 n506__vdd n507__vdd 64.94e-3
rc130 n507__vdd n508__vdd 59.64e-3
rc131 n508__vdd n509__vdd 72.23e-3
rc132 n509__vdd n510__vdd 64.94e-3
rc133 n510__vdd n485__vdd 65.29e-3
rc134 n485__vdd vdd 2.634e-3
rc135 vdd n511__vdd 2.88e-3
rc136 n511__vdd n512__vdd 28.26e-3
rc137 n511__vdd n513__vdd 4.908e-3
rc138 n513__vdd n427__vdd 55.25e-3
rc139 n512__vdd n486__vdd 27.99e-3
rc140 n427__vdd n421__vdd 66.16e-3
rc141 n421__vdd n175__vdd 73.44e-3
rc142 n175__vdd n169__vdd 60.85e-3
rc143 n169__vdd n163__vdd 66.16e-3
rc144 n163__vdd n145__vdd 73.44e-3
rc145 n145__vdd n37__vdd 69.85e-3
rc146 n37__vdd n31__vdd 66.16e-3
rc147 n31__vdd n25__vdd 73.44e-3
rc148 n25__vdd n19__vdd 60.85e-3
rc149 n19__vdd n13__vdd 66.16e-3
rc150 n13__vdd n7__vdd 73.44e-3
rc151 n7__vdd n514__vdd 55.96e-3
rc152 n514__vdd n515__vdd 2.958e-3
rc153 n514__vdd n498__vdd 6.228e-3
rc154 n429__vdd n486__vdd 7.778e-3
rc155 n423__vdd n487__vdd 7.778e-3
rc156 n177__vdd n488__vdd 7.778e-3
rc157 n171__vdd n489__vdd 7.778e-3
rc158 n165__vdd n490__vdd 7.778e-3
rc159 n147__vdd n491__vdd 7.778e-3
rc160 n39__vdd n492__vdd 7.778e-3
rc161 n33__vdd n493__vdd 7.778e-3
rc162 n27__vdd n494__vdd 7.778e-3
rc163 n21__vdd n495__vdd 7.778e-3
rc164 n15__vdd n496__vdd 7.778e-3
rc165 n9__vdd n497__vdd 7.778e-3
rc166 n3__vdd n498__vdd 7.778e-3
rc167 n11__vdd n499__vdd 7.778e-3
rc168 n17__vdd n500__vdd 7.778e-3
rc169 n23__vdd n501__vdd 7.778e-3
rc170 n29__vdd n502__vdd 7.778e-3
rc171 n35__vdd n503__vdd 7.778e-3
rc172 n41__vdd n504__vdd 7.778e-3
rc173 n149__vdd n505__vdd 7.778e-3
rc174 n167__vdd n506__vdd 7.778e-3
rc175 n173__vdd n507__vdd 7.778e-3
rc176 n179__vdd n508__vdd 7.778e-3
rc177 n425__vdd n509__vdd 7.778e-3
rc178 n431__vdd n510__vdd 7.778e-3
rc179 n482__vdd n511__vdd 7.778e-3
rc180 n481__vdd n513__vdd 7.778e-3
rc181 n2__vdd n515__vdd 7.778e-3
rc183 n2111__vddio vddio 4.041e-3
rc186 vddio n2110__vddio 5.514e-3
rc188 n2110__vddio n2116__vddio 65.23e-3
rc189 n2116__vddio n2117__vddio 66.22e-3
rc190 n2117__vddio n2118__vddio 73.5e-3
rc191 n2118__vddio n2119__vddio 60.92e-3
rc192 n2119__vddio n2120__vddio 66.22e-3
rc193 n2120__vddio n2121__vddio 73.5e-3
rc194 n2121__vddio n2122__vddio 69.91e-3
rc195 n2122__vddio n2123__vddio 66.22e-3
rc196 n2123__vddio n2124__vddio 73.5e-3
rc197 n2124__vddio n2125__vddio 60.92e-3
rc198 n2125__vddio n2126__vddio 66.22e-3
rc199 n2126__vddio n2127__vddio 73.5e-3
rc200 n2127__vddio n209__vddio 51.98e-3
rc202 n209__vddio n2129__vddio 5.514e-3
rc204 n2129__vddio vddio 4.908e-3
rc207 n2129__vddio n2133__vddio 49.67e-3
rc208 vddio n2134__vddio 60.94e-3
rc209 n2133__vddio n2135__vddio 73.44e-3
rc210 n2134__vddio n455__vddio 72.72e-3
rc211 n2135__vddio n2136__vddio 66.16e-3
rc212 n455__vddio n2137__vddio 66.88e-3
rc213 n2136__vddio n2138__vddio 60.85e-3
rc214 n2137__vddio n2139__vddio 60.85e-3
rc215 n2138__vddio n2140__vddio 73.44e-3
rc216 n2139__vddio n2141__vddio 73.44e-3
rc217 n2140__vddio n2142__vddio 66.16e-3
rc218 n2141__vddio n2143__vddio 66.16e-3
rc219 n2142__vddio n2144__vddio 69.85e-3
rc220 n2143__vddio n2145__vddio 69.85e-3
rc221 n2144__vddio n2146__vddio 73.44e-3
rc222 n2145__vddio n2147__vddio 73.44e-3
rc223 n2146__vddio n2148__vddio 66.16e-3
rc224 n2147__vddio n2149__vddio 66.16e-3
rc225 n2148__vddio n2150__vddio 60.85e-3
rc226 n2149__vddio n2151__vddio 60.85e-3
rc227 n2150__vddio n2152__vddio 73.44e-3
rc228 n2151__vddio n2153__vddio 73.44e-3
rc229 n2152__vddio n2154__vddio 66.16e-3
rc230 n2153__vddio n2155__vddio 66.16e-3
rc231 n2154__vddio n2156__vddio 28.36e-3
rc232 n2155__vddio n2157__vddio 28.36e-3
rc233 n2156__vddio vddio 24.26e-3
rc234 n2157__vddio n2111__vddio 36.08e-3
rc235 n2105__vddio n2111__vddio 7.778e-3
rc236 n2100__vddio n2111__vddio 7.778e-3
rc237 n2107__vddio vddio 7.778e-3
rc238 n2102__vddio vddio 7.778e-3
rc239 n2104__vddio n2110__vddio 7.778e-3
rc240 n1724__vddio n2116__vddio 7.778e-3
rc241 n1676__vddio n2117__vddio 7.778e-3
rc242 n1407__vddio n2118__vddio 7.778e-3
rc243 n1292__vddio n2119__vddio 7.778e-3
rc244 n1198__vddio n2120__vddio 7.778e-3
rc245 n1030__vddio n2121__vddio 7.778e-3
rc246 n912__vddio n2122__vddio 7.778e-3
rc247 n825__vddio n2123__vddio 7.778e-3
rc248 n647__vddio n2124__vddio 7.778e-3
rc249 n574__vddio n2125__vddio 7.778e-3
rc250 n459__vddio n2126__vddio 7.778e-3
rc251 n281__vddio n2127__vddio 7.778e-3
rc252 n93__vddio n209__vddio 7.778e-3
rc253 n206__vddio n2129__vddio 7.778e-3
rc254 n91__vddio n2129__vddio 7.778e-3
rc255 n204__vddio vddio 7.778e-3
rc256 n89__vddio vddio 7.778e-3
rc257 n279__vddio n2133__vddio 7.778e-3
rc258 n277__vddio n2134__vddio 7.778e-3
rc259 n457__vddio n2135__vddio 7.778e-3
rc260 n572__vddio n2136__vddio 7.778e-3
rc261 n570__vddio n2137__vddio 7.778e-3
rc262 n645__vddio n2138__vddio 7.778e-3
rc263 n643__vddio n2139__vddio 7.778e-3
rc264 n823__vddio n2140__vddio 7.778e-3
rc265 n821__vddio n2141__vddio 7.778e-3
rc266 n910__vddio n2142__vddio 7.778e-3
rc267 n908__vddio n2143__vddio 7.778e-3
rc268 n1028__vddio n2144__vddio 7.778e-3
rc269 n1026__vddio n2145__vddio 7.778e-3
rc270 n1196__vddio n2146__vddio 7.778e-3
rc271 n1194__vddio n2147__vddio 7.778e-3
rc272 n1290__vddio n2148__vddio 7.778e-3
rc273 n1288__vddio n2149__vddio 7.778e-3
rc274 n1405__vddio n2150__vddio 7.778e-3
rc275 n1403__vddio n2151__vddio 7.778e-3
rc276 n1674__vddio n2152__vddio 7.778e-3
rc277 n1672__vddio n2153__vddio 7.778e-3
rc278 n1722__vddio n2154__vddio 7.778e-3
rc279 n1720__vddio n2155__vddio 7.778e-3
rd2 n89__vddio n91__vddio 26.8e-3
rd4 n91__vddio n93__vddio 30.11e-3
rd5 n93__vddio n94__vddio 13.89e-3
rd6 n1__vdd n2__vdd 13.89e-3
rd7 n2__vdd n3__vdd 27.06e-3
rd9 n3__vdd n5__vdd 30.4e-3
rd10 n5__vdd n6__vdd 7.778e-3
rd12 n204__vddio n206__vddio 27.06e-3
rd14 n206__vddio n208__vddio 30.4e-3
rd15 n208__vddio n209__vddio 7.778e-3
rd16 n7__vdd n8__vdd 7.778e-3
rd17 n8__vdd n9__vdd 27.06e-3
rd19 n9__vdd n11__vdd 30.4e-3
rd20 n11__vdd n12__vdd 13.89e-3
rd22 n277__vddio n279__vddio 27.06e-3
rd24 n279__vddio n281__vddio 30.4e-3
rd25 n281__vddio n282__vddio 13.89e-3
rd26 n13__vdd n14__vdd 7.778e-3
rd27 n14__vdd n15__vdd 27.06e-3
rd29 n15__vdd n17__vdd 30.4e-3
rd30 n17__vdd n18__vdd 13.89e-3
rd31 n455__vddio n456__vddio 7.778e-3
rd32 n456__vddio n457__vddio 27.24e-3
rd34 n457__vddio n459__vddio 30.4e-3
rd35 n459__vddio n460__vddio 13.89e-3
rd36 n19__vdd n20__vdd 7.778e-3
rd37 n20__vdd n21__vdd 27.06e-3
rd39 n21__vdd n23__vdd 30.4e-3
rd40 n23__vdd n24__vdd 13.89e-3
rd42 n570__vddio n572__vddio 27.06e-3
rd44 n572__vddio n574__vddio 30.4e-3
rd45 n574__vddio n575__vddio 13.89e-3
rd46 n25__vdd n26__vdd 7.778e-3
rd47 n26__vdd n27__vdd 27.06e-3
rd49 n27__vdd n29__vdd 30.4e-3
rd50 n29__vdd n30__vdd 13.89e-3
rd52 n643__vddio n645__vddio 27.06e-3
rd54 n645__vddio n647__vddio 30.4e-3
rd55 n647__vddio n648__vddio 13.89e-3
rd56 n31__vdd n32__vdd 7.778e-3
rd57 n32__vdd n33__vdd 27.06e-3
rd59 n33__vdd n35__vdd 30.4e-3
rd60 n35__vdd n36__vdd 13.89e-3
rd62 n821__vddio n823__vddio 27.06e-3
rd64 n823__vddio n825__vddio 30.4e-3
rd65 n825__vddio n826__vddio 13.89e-3
rd66 n1537__chipdriverout n1577__chipdriverout 11.67e-3
rd67 n37__vdd n38__vdd 7.778e-3
rd68 n38__vdd n39__vdd 27.06e-3
rd70 n39__vdd n41__vdd 30.4e-3
rd71 n41__vdd n42__vdd 13.89e-3
rd73 n908__vddio n910__vddio 27.06e-3
rd75 n910__vddio n912__vddio 30.4e-3
rd76 n912__vddio n913__vddio 13.89e-3
rd78 n547__vss n549__vss 27.06e-3
rd80 n549__vss n551__vss 30.4e-3
rd81 n551__vss n552__vss 13.89e-3
rd82 n145__vdd n146__vdd 7.778e-3
rd83 n146__vdd n147__vdd 27.06e-3
rd85 n147__vdd n149__vdd 30.4e-3
rd86 n149__vdd n150__vdd 13.89e-3
rd88 n1026__vddio n1028__vddio 27.06e-3
rd90 n1028__vddio n1030__vddio 30.4e-3
rd91 n1030__vddio n1031__vddio 13.89e-3
rd92 n163__vdd n164__vdd 7.778e-3
rd93 n164__vdd n165__vdd 27.06e-3
rd95 n165__vdd n167__vdd 30.4e-3
rd96 n167__vdd n168__vdd 13.89e-3
rd98 n1194__vddio n1196__vddio 27.06e-3
rd100 n1196__vddio n1198__vddio 30.4e-3
rd101 n1198__vddio n1199__vddio 13.89e-3
rd102 n169__vdd n170__vdd 7.778e-3
rd103 n170__vdd n171__vdd 27.06e-3
rd105 n171__vdd n173__vdd 30.4e-3
rd106 n173__vdd n174__vdd 13.89e-3
rd108 n1288__vddio n1290__vddio 27.06e-3
rd110 n1290__vddio n1292__vddio 30.4e-3
rd111 n1292__vddio n1293__vddio 13.89e-3
rd112 n175__vdd n176__vdd 7.778e-3
rd113 n176__vdd n177__vdd 27.06e-3
rd115 n177__vdd n179__vdd 30.4e-3
rd116 n179__vdd n180__vdd 13.89e-3
rd118 n1403__vddio n1405__vddio 27.06e-3
rd120 n1405__vddio n1407__vddio 30.4e-3
rd121 n1407__vddio n1408__vddio 13.89e-3
rd122 n421__vdd n422__vdd 7.778e-3
rd123 n422__vdd n423__vdd 27.06e-3
rd125 n423__vdd n425__vdd 30.4e-3
rd126 n425__vdd n426__vdd 13.89e-3
rd128 n1672__vddio n1674__vddio 27.06e-3
rd130 n1674__vddio n1676__vddio 30.4e-3
rd131 n1676__vddio n1677__vddio 13.89e-3
rd132 n1312__vss n1313__vss 14.16e-3
rd133 n1313__vss n1314__vss 68.49e-3
rd134 n1314__vss n1315__vss 55.79e-3
rd135 n1315__vss n1316__vss 9.752e-3
rd136 n1316__vss n1317__vss 30.4e-3
rd138 n1317__vss n1319__vss 27.06e-3
rd140 n1319__vss n1321__vss 30.4e-3
rd142 n1312__vss n1323__vss 30.4e-3
rd144 n1323__vss n1325__vss 27.06e-3
rd146 n1325__vss n1327__vss 30.4e-3
rd148 n1327__vss n1329__vss 44.29e-3
rd150 n1315__vss n1330__vss 31.42e-3
rd151 n1330__vss n1331__vss 97.75e-3
rd152 n1331__vss n1332__vss 14.16e-3
rd153 n1332__vss n1333__vss 30.4e-3
rd155 n1333__vss n1335__vss 27.06e-3
rd157 n1335__vss n1337__vss 30.4e-3
rd159 n1331__vss n1339__vss 90.2e-3
rd160 n1339__vss n1340__vss 24.82e-3
rd161 n1340__vss n1341__vss 9.752e-3
rd162 n1341__vss n1342__vss 30.4e-3
rd164 n1342__vss n1344__vss 27.06e-3
rd166 n1344__vss n1346__vss 30.4e-3
rd168 n1340__vss n1348__vss 63.55e-3
rd169 n1348__vss n1349__vss 55.75e-3
rd170 n1349__vss n1350__vss 9.793e-3
rd171 n1350__vss n1351__vss 30.4e-3
rd173 n1351__vss n1353__vss 27.06e-3
rd175 n1353__vss n1355__vss 30.4e-3
rd177 n1349__vss n1357__vss 30.67e-3
rd178 n1357__vss n1358__vss 98.59e-3
rd179 n1358__vss n1359__vss 27.52e-3
rd180 n1358__vss n1360__vss 98.59e-3
rd181 n1360__vss n1361__vss 40.08e-3
rd182 n1361__vss n1362__vss 10.97e-3
rd183 n1362__vss n1363__vss 30.4e-3
rd185 n1363__vss n1365__vss 27.06e-3
rd187 n1365__vss n1367__vss 30.4e-3
rd189 n1361__vss n1369__vss 43.11e-3
rd190 n1369__vss n1370__vss 82.62e-3
rd191 n1370__vss n1371__vss 14.45e-3
rd192 n1371__vss n1372__vss 30.4e-3
rd194 n1372__vss n1374__vss 27.06e-3
rd196 n1374__vss n1376__vss 30.4e-3
rd198 n1370__vss n1378__vss 98.59e-3
rd199 n1378__vss n1379__vss 18.46e-3
rd200 n1379__vss n1380__vss 11.75e-3
rd201 n1380__vss n1381__vss 30.4e-3
rd203 n1381__vss n1383__vss 27.06e-3
rd205 n1383__vss n1385__vss 30.4e-3
rd207 n1379__vss n1387__vss 62.82e-3
rd208 n1387__vss n1388__vss 39.29e-3
rd209 n1388__vss n1389__vss 11.86e-3
rd210 n1389__vss n1390__vss 30.4e-3
rd212 n1390__vss n1392__vss 27.06e-3
rd214 n1392__vss n1394__vss 30.4e-3
rd216 n1388__vss n1396__vss 41.7e-3
rd217 n1396__vss n1397__vss 81.09e-3
rd218 n1397__vss n1398__vss 14.01e-3
rd219 n1398__vss n1399__vss 30.4e-3
rd221 n1399__vss n1401__vss 27.06e-3
rd223 n1401__vss n1403__vss 30.4e-3
rd225 n1397__vss n1405__vss 98.59e-3
rd226 n1405__vss n1406__vss 18.95e-3
rd227 n1406__vss n1407__vss 11.63e-3
rd228 n1407__vss n1408__vss 30.4e-3
rd230 n1408__vss n1410__vss 27.06e-3
rd232 n1410__vss n1412__vss 30.4e-3
rd234 n1406__vss n1414__vss 62.61e-3
rd235 n1414__vss n1415__vss 98.12e-3
rd236 n1415__vss n1416__vss 14.16e-3
rd237 n1416__vss n1417__vss 30.4e-3
rd239 n1417__vss n1419__vss 27.06e-3
rd241 n1419__vss n1421__vss 30.4e-3
rd243 n427__vdd n428__vdd 7.778e-3
rd244 n428__vdd n429__vdd 27.06e-3
rd246 n429__vdd n431__vdd 30.4e-3
rd247 n431__vdd n432__vdd 13.89e-3
rd249 n1720__vddio n1722__vddio 27.06e-3
rd251 n1722__vddio n1724__vddio 30.4e-3
rd252 n1724__vddio n1725__vddio 13.89e-3
rd254 n2100__vddio n2102__vddio 27.06e-3
rd256 n2102__vddio n2104__vddio 30.4e-3
rd257 n2104__vddio n2027__vddio 13.89e-3
rd258 n2045__vddio n2100__vddio 13.89e-3
rd259 n2071__vddio n2102__vddio 13.89e-3
rd260 n434__vdd n481__vdd 13.89e-3
rd261 n481__vdd n482__vdd 27.06e-3
rd263 n482__vdd n484__vdd 30.4e-3
rd264 n484__vdd n485__vdd 7.778e-3
rd265 n462__vdd n482__vdd 13.89e-3
rd266 n478__vdd n484__vdd 13.89e-3
rd268 n2016__vss n2018__vss 109.7e-3
rd269 n2018__vss n2019__vss 4.667e-3
rd270 n1928__vss n2016__vss 8.333e-3
rd271 n2002__vss n2018__vss 8.333e-3
rd272 n1861__vss n2020__vss 44.29e-3
rd274 n2020__vss n2001__vss 27.06e-3
rd276 n2001__vss n2023__vss 30.4e-3
rd278 n2023__vss n2009__vss 44.29e-3
rd280 n2009__vss n2026__vss 21.08e-3
rd282 n2026__vss n2028__vss 63.41e-3
rd284 n2028__vss n2015__vss 83.47e-3
rd286 n2015__vss n2031__vss 21.29e-3
rd288 n2031__vss n2033__vss 44.29e-3
rd290 n2033__vss n2035__vss 30.4e-3
rd292 n2035__vss n2037__vss 27.06e-3
rd294 n2037__vss n1863__vss 44.29e-3
rd295 n1925__vss n2020__vss 13.89e-3
rd296 n2007__vss n2023__vss 13.89e-3
rd297 n2011__vss n2026__vss 16.67e-3
rd298 n2013__vss n2028__vss 8.333e-3
rd299 n2005__vss n2031__vss 13.89e-3
rd300 n1931__vss n2033__vss 13.89e-3
rd301 n1973__vss n2035__vss 13.89e-3
rd302 n1946__vss n2037__vss 13.89e-3
rd304 n2105__vddio n2107__vddio 27.06e-3
rd306 n2107__vddio n2109__vddio 30.4e-3
rd307 n2109__vddio n2110__vddio 7.778e-3
rd308 n2043__vddio n2105__vddio 13.89e-3
rd309 n2069__vddio n2107__vddio 13.89e-3
rd310 n2025__vddio n2109__vddio 13.89e-3
re1 n1497__chipdriverout n1537__chipdriverout 20.83e-3
re3 n1861__vss n1863__vss 194.4e-3
re5 n1863__vss n1865__vss 224.7e-3
re7 n1865__vss n1867__vss 4.917e-3
re9 n1867__vss n1869__vss 66.3e-3
re11 n1869__vss n1871__vss 59.18e-3
re13 n1871__vss n1873__vss 35.78e-3
re15 n1873__vss n1875__vss 94.95e-3
re17 n1875__vss n1877__vss 8.478e-3
re19 n1877__vss n1879__vss 86.47e-3
re21 n1879__vss n1881__vss 28.99e-3
re23 n1881__vss n1883__vss 65.96e-3
re25 n1883__vss n1885__vss 59.51e-3
re27 n1885__vss n1887__vss 35.44e-3
re29 n1887__vss n1889__vss 94.95e-3
re31 n1889__vss n1359__vss 8.817e-3
re33 n1359__vss n1892__vss 86.13e-3
re35 n1892__vss n1894__vss 46.29e-3
re37 n1894__vss n1896__vss 48.66e-3
re39 n1896__vss n1898__vss 76.81e-3
re41 n1898__vss n1900__vss 18.14e-3
re43 n1900__vss n1902__vss 94.95e-3
re45 n1902__vss n1904__vss 26.11e-3
re47 n1904__vss n1906__vss 68.84e-3
re49 n1906__vss n1908__vss 46.63e-3
re51 n1908__vss n1910__vss 48.32e-3
re53 n1910__vss n1912__vss 77.15e-3
re55 n1912__vss n1914__vss 17.8e-3
re57 n1914__vss n1916__vss 94.95e-3
re59 n1916__vss n1918__vss 26.45e-3
re61 n1918__vss n1920__vss 68.5e-3
re63 n1920__vss n1922__vss 94.95e-3
re65 n1922__vss n1924__vss 6.782e-3
re66 n1924__vss n1416__vss 13.89e-3
re67 n1817__vss n1861__vss 13.89e-3
re68 n1839__vss n1863__vss 13.89e-3
re69 n1461__vss n1865__vss 16.67e-3
re70 n1313__vss n1865__vss 16.67e-3
re71 n1312__vss n1867__vss 13.89e-3
re72 n1459__vss n1867__vss 13.89e-3
re73 n1471__vss n1869__vss 8.333e-3
re74 n1314__vss n1869__vss 8.333e-3
re75 n1473__vss n1871__vss 13.89e-3
re76 n1316__vss n1871__vss 13.89e-3
re77 n1330__vss n1873__vss 8.333e-3
re78 n1477__vss n1873__vss 8.333e-3
re79 n1479__vss n1875__vss 8.333e-3
re80 n1331__vss n1875__vss 8.333e-3
re81 n1481__vss n1877__vss 13.89e-3
re82 n1332__vss n1877__vss 13.89e-3
re83 n1339__vss n1879__vss 8.333e-3
re84 n1485__vss n1879__vss 8.333e-3
re85 n1341__vss n1881__vss 13.89e-3
re86 n1487__vss n1881__vss 13.89e-3
re87 n1491__vss n1883__vss 8.333e-3
re88 n1348__vss n1883__vss 8.333e-3
re89 n1493__vss n1885__vss 13.89e-3
re90 n1350__vss n1885__vss 13.89e-3
re91 n1357__vss n1887__vss 8.333e-3
re92 n1497__vss n1887__vss 8.333e-3
re93 n1499__vss n1889__vss 8.333e-3
re94 n1358__vss n1889__vss 8.333e-3
re95 n1501__vss n1359__vss 13.89e-3
re96 n1505__vss n1892__vss 8.333e-3
re97 n1360__vss n1892__vss 8.333e-3
re98 n1507__vss n1894__vss 13.89e-3
re99 n1362__vss n1894__vss 13.89e-3
re100 n1511__vss n1896__vss 8.333e-3
re101 n1369__vss n1896__vss 8.333e-3
re102 n1513__vss n1898__vss 13.89e-3
re103 n1371__vss n1898__vss 13.89e-3
re104 n1370__vss n1900__vss 8.333e-3
re105 n1514__vss n1900__vss 8.333e-3
re106 n1519__vss n1902__vss 8.333e-3
re107 n1378__vss n1902__vss 8.333e-3
re108 n1521__vss n1904__vss 13.89e-3
re109 n1380__vss n1904__vss 13.89e-3
re110 n1525__vss n1906__vss 8.333e-3
re111 n1387__vss n1906__vss 8.333e-3
re112 n1527__vss n1908__vss 13.89e-3
re113 n1389__vss n1908__vss 13.89e-3
re114 n1531__vss n1910__vss 8.333e-3
re115 n1396__vss n1910__vss 8.333e-3
re116 n1533__vss n1912__vss 13.89e-3
re117 n1398__vss n1912__vss 13.89e-3
re118 n1397__vss n1914__vss 8.333e-3
re119 n1534__vss n1914__vss 8.333e-3
re120 n1539__vss n1916__vss 8.333e-3
re121 n1405__vss n1916__vss 8.333e-3
re122 n1541__vss n1918__vss 13.89e-3
re123 n1407__vss n1918__vss 13.89e-3
re124 n1414__vss n1920__vss 8.333e-3
re125 n1545__vss n1920__vss 8.333e-3
re126 n1415__vss n1922__vss 8.333e-3
re127 n1547__vss n1922__vss 8.333e-3
re128 n1549__vss n1924__vss 13.89e-3
re130 n1925__vss n1927__vss 66.75e-3
re131 n1927__vss n1928__vss 84.47e-3
re133 n1928__vss n1930__vss 160.8e-3
re134 n1930__vss n1931__vss 126.1e-3
re136 n1931__vss n1933__vss 242.8e-3
re138 n1933__vss n1476__vss 186.7e-3
re140 n1476__vss n1484__vss 207.3e-3
re142 n1484__vss n1490__vss 171.7e-3
re144 n1490__vss n1496__vss 186.7e-3
re146 n1496__vss n552__vss 207.3e-3
re148 n552__vss n1510__vss 197.1e-3
re150 n1510__vss n1518__vss 186.7e-3
re152 n1518__vss n1524__vss 207.3e-3
re154 n1524__vss n1530__vss 171.7e-3
re156 n1530__vss n1538__vss 186.7e-3
re158 n1538__vss n1544__vss 207.3e-3
re160 n1544__vss n1552__vss 253.7e-3
re162 n1927__vss n1946__vss 126.6e-3
re164 n1946__vss n1948__vss 242.9e-3
re166 n1948__vss n1950__vss 186.8e-3
re168 n1950__vss n1952__vss 207.4e-3
re170 n1952__vss n1954__vss 171.8e-3
re172 n1954__vss n1956__vss 186.8e-3
re174 n1956__vss n1958__vss 207.4e-3
re176 n1958__vss n1960__vss 197.2e-3
re178 n1960__vss n1962__vss 186.8e-3
re180 n1962__vss n1964__vss 207.4e-3
re182 n1964__vss n1966__vss 171.8e-3
re184 n1966__vss n1968__vss 186.8e-3
re186 n1968__vss n1970__vss 207.4e-3
re188 n1970__vss n1972__vss 253.8e-3
re189 n1972__vss n1417__vss 13.89e-3
re190 n1928__vss n1973__vss 127.2e-3
re192 n1973__vss n1975__vss 243.1e-3
re194 n1975__vss n1977__vss 187e-3
re196 n1977__vss n1979__vss 207.5e-3
re198 n1979__vss n1981__vss 172e-3
re200 n1981__vss n1983__vss 187e-3
re202 n1983__vss n1985__vss 207.5e-3
re204 n1985__vss n1987__vss 197.4e-3
re206 n1987__vss n1989__vss 187e-3
re208 n1989__vss n1991__vss 207.5e-3
re210 n1991__vss n1993__vss 172e-3
re212 n1993__vss n1995__vss 187e-3
re214 n1995__vss n1997__vss 207.5e-3
re216 n1997__vss n1999__vss 254e-3
re217 n1999__vss n1419__vss 13.89e-3
re218 n1928__vss n2000__vss 67.35e-3
re219 n2000__vss n2001__vss 13.89e-3
re220 n1930__vss n2002__vss 90.18e-3
re222 n2002__vss n2004__vss 138.7e-3
re223 n2004__vss n2005__vss 126.6e-3
re225 n1930__vss n2007__vss 66.16e-3
re226 n2007__vss n1831__vss 13.89e-3
re227 n2004__vss n2008__vss 66.68e-3
re228 n2008__vss n2009__vss 13.89e-3
re229 n2005__vss n1470__vss 242.8e-3
re231 n1818__vss n1925__vss 13.89e-3
re232 n1848__vss n1928__vss 8.333e-3
re233 n1845__vss n1931__vss 13.89e-3
re234 n1327__vss n1933__vss 13.89e-3
re235 n1467__vss n1933__vss 13.89e-3
re236 n1321__vss n1476__vss 13.89e-3
re237 n1337__vss n1484__vss 13.89e-3
re238 n1346__vss n1490__vss 13.89e-3
re239 n1355__vss n1496__vss 13.89e-3
re240 n1367__vss n1510__vss 13.89e-3
re241 n1376__vss n1518__vss 13.89e-3
re242 n1385__vss n1524__vss 13.89e-3
re243 n1394__vss n1530__vss 13.89e-3
re244 n1403__vss n1538__vss 13.89e-3
re245 n1412__vss n1544__vss 13.89e-3
re246 n1421__vss n1552__vss 13.89e-3
re247 n1841__vss n1946__vss 13.89e-3
re248 n1463__vss n1948__vss 13.89e-3
re249 n1323__vss n1948__vss 13.89e-3
re250 n1317__vss n1950__vss 13.89e-3
re251 n1474__vss n1950__vss 13.89e-3
re252 n1482__vss n1952__vss 13.89e-3
re253 n1333__vss n1952__vss 13.89e-3
re254 n1488__vss n1954__vss 13.89e-3
re255 n1342__vss n1954__vss 13.89e-3
re256 n1351__vss n1956__vss 13.89e-3
re257 n1494__vss n1956__vss 13.89e-3
re258 n547__vss n1958__vss 13.89e-3
re259 n1502__vss n1958__vss 13.89e-3
re260 n1363__vss n1960__vss 13.89e-3
re261 n1508__vss n1960__vss 13.89e-3
re262 n1516__vss n1962__vss 13.89e-3
re263 n1372__vss n1962__vss 13.89e-3
re264 n1522__vss n1964__vss 13.89e-3
re265 n1381__vss n1964__vss 13.89e-3
re266 n1528__vss n1966__vss 13.89e-3
re267 n1390__vss n1966__vss 13.89e-3
re268 n1399__vss n1968__vss 13.89e-3
re269 n1536__vss n1968__vss 13.89e-3
re270 n1408__vss n1970__vss 13.89e-3
re271 n1542__vss n1970__vss 13.89e-3
re272 n1550__vss n1972__vss 13.89e-3
re273 n1843__vss n1973__vss 13.89e-3
re274 n1325__vss n1975__vss 13.89e-3
re275 n1465__vss n1975__vss 13.89e-3
re276 n1319__vss n1977__vss 13.89e-3
re277 n1475__vss n1977__vss 13.89e-3
re278 n1335__vss n1979__vss 13.89e-3
re279 n1483__vss n1979__vss 13.89e-3
re280 n1489__vss n1981__vss 13.89e-3
re281 n1344__vss n1981__vss 13.89e-3
re282 n1353__vss n1983__vss 13.89e-3
re283 n1495__vss n1983__vss 13.89e-3
re284 n1503__vss n1985__vss 13.89e-3
re285 n549__vss n1985__vss 13.89e-3
re286 n1509__vss n1987__vss 13.89e-3
re287 n1365__vss n1987__vss 13.89e-3
re288 n1374__vss n1989__vss 13.89e-3
re289 n1517__vss n1989__vss 13.89e-3
re290 n1523__vss n1991__vss 13.89e-3
re291 n1383__vss n1991__vss 13.89e-3
re292 n1392__vss n1993__vss 13.89e-3
re293 n1529__vss n1993__vss 13.89e-3
re294 n1401__vss n1995__vss 13.89e-3
re295 n1537__vss n1995__vss 13.89e-3
re296 n1410__vss n1997__vss 13.89e-3
re297 n1543__vss n1997__vss 13.89e-3
re298 n1551__vss n1999__vss 13.89e-3
re299 n1829__vss n2000__vss 13.89e-3
re300 n1850__vss n2002__vss 8.333e-3
re301 n1847__vss n2005__vss 13.89e-3
re302 n1832__vss n2008__vss 13.89e-3
re303 n1329__vss n1470__vss 13.89e-3
re305 n434__vdd n435__vdd 232.7e-3
re306 n435__vdd n436__vdd 186.7e-3
re307 n436__vdd n437__vdd 79.91e-3
re308 n437__vdd n438__vdd 127.4e-3
re309 n438__vdd n439__vdd 13.82e-3
re310 n439__vdd n440__vdd 142.1e-3
re311 n440__vdd n441__vdd 16.04e-3
re312 n441__vdd n442__vdd 125.1e-3
re313 n442__vdd n443__vdd 61.64e-3
re314 n443__vdd n444__vdd 79.4e-3
re315 n444__vdd n445__vdd 127.9e-3
re316 n445__vdd n446__vdd 163.4e-3
re317 n446__vdd n447__vdd 33.72e-3
re318 n447__vdd n448__vdd 107.3e-3
re319 n448__vdd n449__vdd 79.4e-3
re320 n449__vdd n450__vdd 61.64e-3
re321 n450__vdd n451__vdd 141.7e-3
re322 n451__vdd n452__vdd 3.949e-3
re323 n452__vdd n453__vdd 137.5e-3
re324 n453__vdd n454__vdd 34.23e-3
re325 n454__vdd n455__vdd 106.8e-3
re326 n455__vdd n456__vdd 79.91e-3
re327 n456__vdd n457__vdd 61.13e-3
re328 n457__vdd n458__vdd 141.7e-3
re329 n458__vdd n459__vdd 4.443e-3
re330 n459__vdd n460__vdd 137e-3
re331 n460__vdd n1__vdd 86.51e-3
re332 n1__vdd n144__vdd 54.53e-3
re333 n428__vdd n435__vdd 13.89e-3
re334 n422__vdd n436__vdd 13.89e-3
re335 n412__vdd n437__vdd 12.5e-3
re336 n176__vdd n438__vdd 13.89e-3
re337 n414__vdd n439__vdd 12.5e-3
re338 n416__vdd n440__vdd 12.5e-3
re339 n170__vdd n441__vdd 13.89e-3
re340 n418__vdd n442__vdd 12.5e-3
re341 n164__vdd n443__vdd 13.89e-3
re342 n420__vdd n444__vdd 12.5e-3
re343 n146__vdd n445__vdd 13.89e-3
re344 n125__vdd n446__vdd 12.5e-3
re345 n38__vdd n447__vdd 13.89e-3
re346 n127__vdd n448__vdd 12.5e-3
re347 n32__vdd n449__vdd 13.89e-3
re348 n129__vdd n450__vdd 12.5e-3
re349 n131__vdd n451__vdd 12.5e-3
re350 n26__vdd n452__vdd 13.89e-3
re351 n133__vdd n453__vdd 12.5e-3
re352 n20__vdd n454__vdd 13.89e-3
re353 n135__vdd n455__vdd 12.5e-3
re354 n14__vdd n456__vdd 13.89e-3
re355 n137__vdd n457__vdd 12.5e-3
re356 n139__vdd n458__vdd 12.5e-3
re357 n8__vdd n459__vdd 13.89e-3
re358 n141__vdd n460__vdd 12.5e-3
re360 n462__vdd n463__vdd 232.5e-3
re361 n463__vdd n464__vdd 186.5e-3
re362 n464__vdd n465__vdd 207.1e-3
re363 n465__vdd n466__vdd 171.6e-3
re364 n466__vdd n467__vdd 186.5e-3
re365 n467__vdd n468__vdd 207.1e-3
re366 n468__vdd n469__vdd 196.9e-3
re367 n469__vdd n470__vdd 186.5e-3
re368 n470__vdd n471__vdd 207.1e-3
re369 n471__vdd n472__vdd 171.6e-3
re370 n472__vdd n473__vdd 186.5e-3
re371 n473__vdd n474__vdd 207.1e-3
re372 n474__vdd n475__vdd 223.3e-3
re374 n429__vdd n463__vdd 13.89e-3
re375 n423__vdd n464__vdd 13.89e-3
re376 n177__vdd n465__vdd 13.89e-3
re377 n171__vdd n466__vdd 13.89e-3
re378 n165__vdd n467__vdd 13.89e-3
re379 n147__vdd n468__vdd 13.89e-3
re380 n39__vdd n469__vdd 13.89e-3
re381 n33__vdd n470__vdd 13.89e-3
re382 n27__vdd n471__vdd 13.89e-3
re383 n21__vdd n472__vdd 13.89e-3
re384 n15__vdd n473__vdd 13.89e-3
re385 n9__vdd n474__vdd 13.89e-3
re386 n3__vdd n475__vdd 13.89e-3
re388 n478__vdd n432__vdd 231.5e-3
re389 n432__vdd n426__vdd 185.5e-3
re390 n426__vdd n180__vdd 206.1e-3
re391 n180__vdd n174__vdd 170.6e-3
re392 n174__vdd n168__vdd 185.5e-3
re393 n168__vdd n150__vdd 206.1e-3
re394 n150__vdd n42__vdd 195.9e-3
re395 n42__vdd n36__vdd 185.5e-3
re396 n36__vdd n30__vdd 206.1e-3
re397 n30__vdd n24__vdd 170.6e-3
re398 n24__vdd n18__vdd 185.5e-3
re399 n18__vdd n12__vdd 206.1e-3
re400 n12__vdd n479__vdd 222.3e-3
re402 n5__vdd n479__vdd 13.89e-3
re404 n2025__vddio n2027__vddio 187.4e-3
re406 n2027__vddio n1725__vddio 187.1e-3
re408 n1725__vddio n1677__vddio 187.3e-3
re410 n1677__vddio n1408__vddio 208e-3
re412 n1408__vddio n1293__vddio 172.3e-3
re414 n1293__vddio n1199__vddio 187.3e-3
re416 n1199__vddio n1031__vddio 208e-3
re418 n1031__vddio n913__vddio 197.8e-3
re420 n913__vddio n826__vddio 187.3e-3
re422 n826__vddio n648__vddio 208e-3
re424 n648__vddio n575__vddio 172.3e-3
re426 n575__vddio n460__vddio 187.3e-3
re428 n460__vddio n282__vddio 208e-3
re430 n282__vddio n2041__vddio 173.8e-3
re432 n2041__vddio n94__vddio 207.4e-3
re433 n94__vddio n66__vddio 13.89e-3
re434 n2021__vddio n2025__vddio 13.89e-3
re435 n2017__vddio n2027__vddio 13.89e-3
re436 n1726__vddio n1725__vddio 13.89e-3
re437 n1668__vddio n1677__vddio 13.89e-3
re438 n1399__vddio n1408__vddio 13.89e-3
re439 n1286__vddio n1293__vddio 13.89e-3
re440 n1169__vddio n1199__vddio 13.89e-3
re441 n1032__vddio n1031__vddio 13.89e-3
re442 n904__vddio n913__vddio 13.89e-3
re443 n798__vddio n826__vddio 13.89e-3
re444 n639__vddio n648__vddio 13.89e-3
re445 n568__vddio n575__vddio 13.89e-3
re446 n423__vddio n460__vddio 13.89e-3
re447 n273__vddio n282__vddio 13.89e-3
re448 n208__vddio n2041__vddio 13.89e-3
re449 n202__vddio n2041__vddio 13.89e-3
re451 n2043__vddio n2045__vddio 186.7e-3
re453 n2045__vddio n2047__vddio 186.5e-3
re455 n2047__vddio n2049__vddio 186.7e-3
re457 n2049__vddio n2051__vddio 207.3e-3
re459 n2051__vddio n1284__vddio 171.7e-3
re461 n1284__vddio n2054__vddio 186.7e-3
re463 n2054__vddio n2056__vddio 207.3e-3
re465 n2056__vddio n2058__vddio 197.1e-3
re467 n2058__vddio n796__vddio 186.7e-3
re469 n796__vddio n2061__vddio 207.3e-3
re471 n2061__vddio n566__vddio 171.7e-3
re473 n566__vddio n426__vddio 188.9e-3
re475 n426__vddio n2065__vddio 205.4e-3
re477 n2065__vddio n200__vddio 173.3e-3
re479 n200__vddio n64__vddio 206.5e-3
re481 n2024__vddio n2043__vddio 13.89e-3
re482 n2020__vddio n2045__vddio 13.89e-3
re483 n1729__vddio n2047__vddio 13.89e-3
re484 n1720__vddio n2047__vddio 13.89e-3
re485 n1671__vddio n2049__vddio 13.89e-3
re486 n1672__vddio n2049__vddio 13.89e-3
re487 n1403__vddio n2051__vddio 13.89e-3
re488 n1402__vddio n2051__vddio 13.89e-3
re489 n1288__vddio n1284__vddio 13.89e-3
re490 n1172__vddio n2054__vddio 13.89e-3
re491 n1194__vddio n2054__vddio 13.89e-3
re492 n1035__vddio n2056__vddio 13.89e-3
re493 n1026__vddio n2056__vddio 13.89e-3
re494 n908__vddio n2058__vddio 13.89e-3
re495 n907__vddio n2058__vddio 13.89e-3
re496 n821__vddio n796__vddio 13.89e-3
re497 n643__vddio n2061__vddio 13.89e-3
re498 n642__vddio n2061__vddio 13.89e-3
re499 n570__vddio n566__vddio 13.89e-3
re500 n456__vddio n426__vddio 13.89e-3
re501 n277__vddio n2065__vddio 13.89e-3
re502 n276__vddio n2065__vddio 13.89e-3
re503 n204__vddio n200__vddio 13.89e-3
re504 n89__vddio n64__vddio 13.89e-3
re506 n2069__vddio n2071__vddio 186.7e-3
re508 n2071__vddio n2073__vddio 186.5e-3
re510 n2073__vddio n2075__vddio 186.7e-3
re512 n2075__vddio n2077__vddio 207.3e-3
re514 n2077__vddio n2079__vddio 171.7e-3
re516 n2079__vddio n2081__vddio 186.7e-3
re518 n2081__vddio n2083__vddio 207.3e-3
re520 n2083__vddio n2085__vddio 197.1e-3
re522 n2085__vddio n2087__vddio 186.7e-3
re524 n2087__vddio n2089__vddio 207.3e-3
re526 n2089__vddio n2091__vddio 171.7e-3
re528 n2091__vddio n2093__vddio 186.7e-3
re530 n2093__vddio n2095__vddio 207.3e-3
re532 n2095__vddio n2097__vddio 173.3e-3
re534 n2097__vddio n2099__vddio 206.5e-3
re535 n2099__vddio n91__vddio 13.89e-3
re536 n2023__vddio n2069__vddio 13.89e-3
re537 n2019__vddio n2071__vddio 13.89e-3
re538 n1722__vddio n2073__vddio 13.89e-3
re539 n1728__vddio n2073__vddio 13.89e-3
re540 n1674__vddio n2075__vddio 13.89e-3
re541 n1670__vddio n2075__vddio 13.89e-3
re542 n1401__vddio n2077__vddio 13.89e-3
re543 n1405__vddio n2077__vddio 13.89e-3
re544 n1285__vddio n2079__vddio 13.89e-3
re545 n1290__vddio n2079__vddio 13.89e-3
re546 n1196__vddio n2081__vddio 13.89e-3
re547 n1171__vddio n2081__vddio 13.89e-3
re548 n1028__vddio n2083__vddio 13.89e-3
re549 n1034__vddio n2083__vddio 13.89e-3
re550 n906__vddio n2085__vddio 13.89e-3
re551 n910__vddio n2085__vddio 13.89e-3
re552 n823__vddio n2087__vddio 13.89e-3
re553 n797__vddio n2087__vddio 13.89e-3
re554 n641__vddio n2089__vddio 13.89e-3
re555 n645__vddio n2089__vddio 13.89e-3
re556 n567__vddio n2091__vddio 13.89e-3
re557 n572__vddio n2091__vddio 13.89e-3
re558 n425__vddio n2093__vddio 13.89e-3
re559 n457__vddio n2093__vddio 13.89e-3
re560 n275__vddio n2095__vddio 13.89e-3
re561 n279__vddio n2095__vddio 13.89e-3
re562 n201__vddio n2097__vddio 13.89e-3
re563 n206__vddio n2097__vddio 13.89e-3
re564 n65__vddio n2099__vddio 13.89e-3
re566 n2011__vss n2013__vss 212.2e-3
re568 n2013__vss n1860__vss 282.9e-3
re569 n1860__vss n2015__vss 8.333e-3
re570 n1856__vss n2011__vss 16.67e-3
re571 n1858__vss n2013__vss 8.333e-3
rf1 n64__vddio n65__vddio 107.9e-3
rf2 n65__vddio n66__vddio 105.6e-3
rf3 n66__vddio n67__vddio 13.89e-3
rf4 n200__vddio n201__vddio 107.9e-3
rf5 n201__vddio n202__vddio 105.6e-3
rf6 n202__vddio n203__vddio 13.89e-3
rf8 n273__vddio n275__vddio 105.6e-3
rf9 n275__vddio n276__vddio 94.02e-3
rf11 n423__vddio n425__vddio 103.6e-3
rf12 n425__vddio n426__vddio 107.6e-3
rf13 n566__vddio n567__vddio 106.9e-3
rf14 n567__vddio n568__vddio 104.6e-3
rf17 n639__vddio n641__vddio 104.9e-3
rf18 n641__vddio n642__vddio 93.33e-3
rf19 n796__vddio n797__vddio 107.9e-3
rf20 n797__vddio n798__vddio 105.6e-3
rf21 n798__vddio n799__vddio 13.89e-3
rf22 n1497__chipdriverout n1444__chipdriverout 20.83e-3
rf24 n904__vddio n906__vddio 106.2e-3
rf25 n906__vddio n907__vddio 94.55e-3
rf27 n125__vdd n127__vdd 435.8e-3
rf29 n127__vdd n129__vdd 435.8e-3
rf31 n129__vdd n131__vdd 435.8e-3
rf33 n131__vdd n133__vdd 435.8e-3
rf35 n133__vdd n135__vdd 435.8e-3
rf37 n135__vdd n137__vdd 435.8e-3
rf39 n137__vdd n139__vdd 435.8e-3
rf41 n139__vdd n141__vdd 435.8e-3
rf43 n141__vdd n143__vdd 435.8e-3
rf44 n143__vdd n144__vdd 12.5e-3
rf45 n106__vdd n125__vdd 12.5e-3
rf46 n108__vdd n127__vdd 12.5e-3
rf47 n110__vdd n129__vdd 12.5e-3
rf48 n112__vdd n131__vdd 12.5e-3
rf49 n114__vdd n133__vdd 12.5e-3
rf50 n116__vdd n135__vdd 12.5e-3
rf51 n118__vdd n137__vdd 12.5e-3
rf52 n120__vdd n139__vdd 12.5e-3
rf53 n122__vdd n141__vdd 12.5e-3
rf54 n105__vdd n143__vdd 12.5e-3
rf56 n1032__vddio n1034__vddio 105.6e-3
rf57 n1034__vddio n1035__vddio 94.02e-3
rf58 n2__i5__r2 n14__i5__r2 1.2439
rf60 n15__i5__r1 n9__i5__r1 1.2089
rf62 n1169__vddio n1171__vddio 105.6e-3
rf63 n1171__vddio n1172__vddio 94.02e-3
rf64 n1284__vddio n1285__vddio 103.6e-3
rf65 n1285__vddio n1286__vddio 100.9e-3
rf67 n17__i5__r0 n3__i5__r0 3.3264
rf69 n1399__vddio n1401__vddio 105.6e-3
rf70 n1401__vddio n1402__vddio 94.02e-3
rf72 n412__vdd n414__vdd 435.8e-3
rf74 n414__vdd n416__vdd 435.8e-3
rf76 n416__vdd n418__vdd 435.8e-3
rf78 n418__vdd n420__vdd 435.8e-3
rf79 n420__vdd n411__vdd 12.5e-3
rf80 n403__vdd n412__vdd 12.5e-3
rf81 n405__vdd n414__vdd 12.5e-3
rf82 n407__vdd n416__vdd 12.5e-3
rf83 n409__vdd n418__vdd 12.5e-3
rf85 n1668__vddio n1670__vddio 105.6e-3
rf86 n1670__vddio n1671__vddio 94.02e-3
rf88 n1459__vss n1461__vss 33.06e-3
rf90 n1459__vss n1463__vss 105.6e-3
rf92 n1463__vss n1465__vss 94.02e-3
rf94 n1465__vss n1467__vss 105.6e-3
rf96 n1467__vss n1469__vss 153.9e-3
rf97 n1469__vss n1470__vss 13.89e-3
rf98 n1459__vss n1471__vss 145e-3
rf100 n1471__vss n1473__vss 129.4e-3
rf101 n1473__vss n1474__vss 105.6e-3
rf102 n1474__vss n1475__vss 94.02e-3
rf103 n1475__vss n1476__vss 119.5e-3
rf104 n1473__vss n1477__vss 78.24e-3
rf106 n1477__vss n1479__vss 207.6e-3
rf108 n1479__vss n1481__vss 18.54e-3
rf109 n1481__vss n1482__vss 105.6e-3
rf110 n1482__vss n1483__vss 94.02e-3
rf111 n1483__vss n1484__vss 119.5e-3
rf112 n1481__vss n1485__vss 189.1e-3
rf114 n1485__vss n1487__vss 62.95e-3
rf115 n1487__vss n1488__vss 90.57e-3
rf116 n1488__vss n1489__vss 93.01e-3
rf117 n1489__vss n1490__vss 118.5e-3
rf118 n1487__vss n1491__vss 145.2e-3
rf120 n1491__vss n1493__vss 130.2e-3
rf121 n1493__vss n1494__vss 105.6e-3
rf122 n1494__vss n1495__vss 94.02e-3
rf123 n1495__vss n1496__vss 119.5e-3
rf124 n1493__vss n1497__vss 77.5e-3
rf126 n1497__vss n1499__vss 207.6e-3
rf128 n1499__vss n1501__vss 19.28e-3
rf129 n1501__vss n1502__vss 104.9e-3
rf130 n1502__vss n1503__vss 93.33e-3
rf131 n1503__vss n552__vss 118.8e-3
rf132 n1501__vss n1505__vss 188.4e-3
rf134 n1505__vss n1507__vss 101.2e-3
rf135 n1507__vss n1508__vss 105.6e-3
rf136 n1508__vss n1509__vss 94.02e-3
rf137 n1509__vss n1510__vss 119.5e-3
rf138 n1507__vss n1511__vss 106.4e-3
rf140 n1511__vss n1513__vss 167.5e-3
rf141 n1513__vss n1514__vss 18.18e-3
rf143 n1513__vss n1516__vss 90.57e-3
rf144 n1516__vss n1517__vss 93.01e-3
rf145 n1517__vss n1518__vss 118.5e-3
rf146 n1514__vss n1519__vss 207.6e-3
rf148 n1519__vss n1521__vss 58.05e-3
rf149 n1521__vss n1522__vss 90.57e-3
rf150 n1522__vss n1523__vss 93.01e-3
rf151 n1523__vss n1524__vss 118.5e-3
rf152 n1521__vss n1525__vss 150.1e-3
rf154 n1525__vss n1527__vss 102e-3
rf155 n1527__vss n1528__vss 105.6e-3
rf156 n1528__vss n1529__vss 94.02e-3
rf157 n1529__vss n1530__vss 119.5e-3
rf158 n1527__vss n1531__vss 105.7e-3
rf160 n1531__vss n1533__vss 168.7e-3
rf161 n1533__vss n1534__vss 38.93e-3
rf163 n1533__vss n1536__vss 104.9e-3
rf164 n1536__vss n1537__vss 93.33e-3
rf165 n1537__vss n1538__vss 118.8e-3
rf166 n1534__vss n1539__vss 207.6e-3
rf168 n1539__vss n1541__vss 57.84e-3
rf169 n1541__vss n1542__vss 105.6e-3
rf170 n1542__vss n1543__vss 94.02e-3
rf171 n1543__vss n1544__vss 119.5e-3
rf172 n1541__vss n1545__vss 149.8e-3
rf174 n1545__vss n1547__vss 207.6e-3
rf176 n1547__vss n1549__vss 25.96e-3
rf177 n1549__vss n1550__vss 105.6e-3
rf178 n1550__vss n1551__vss 94.02e-3
rf179 n1551__vss n1552__vss 119.5e-3
rf181 n1726__vddio n1728__vddio 106.2e-3
rf182 n1728__vddio n1729__vddio 94.55e-3
rf184 n1839__vss n1841__vss 104.9e-3
rf186 n1841__vss n1843__vss 93.33e-3
rf188 n1843__vss n1845__vss 104.9e-3
rf190 n1845__vss n1847__vss 153.2e-3
rf191 n1847__vss n1827__vss 13.89e-3
rf192 n1816__vss n1839__vss 13.89e-3
rf193 n1822__vss n1841__vss 13.89e-3
rf194 n1828__vss n1843__vss 13.89e-3
rf195 n1830__vss n1845__vss 13.89e-3
rf197 n2017__vddio n2019__vddio 105.6e-3
rf198 n2019__vddio n2020__vddio 94.02e-3
rf199 n1986__vddio n2017__vddio 13.89e-3
rf201 n1848__vss n1850__vss 307.7e-3
rf202 n1850__vss n1824__vss 8.333e-3
rf203 n1820__vss n1848__vss 8.333e-3
rf205 n1817__vss n1818__vss 104.3e-3
rf207 n1818__vss n1829__vss 92.7e-3
rf209 n1829__vss n1831__vss 104.3e-3
rf211 n1831__vss n1832__vss 152.6e-3
rf214 n1856__vss n1858__vss 207.9e-3
rf216 n1858__vss n1838__vss 277.2e-3
rf217 n1838__vss n1860__vss 8.333e-3
rf218 n1833__vss n1856__vss 16.67e-3
rf219 n1835__vss n1858__vss 8.333e-3
rf221 n2021__vddio n2023__vddio 105.6e-3
rf222 n2023__vddio n2024__vddio 94.02e-3
rf223 n1983__vddio n2021__vddio 13.89e-3
rg1 n1443__chipdriverout n1444__chipdriverout 41.67e-3
rg2 n2__i5__r0 n3__i5__r0 125e-3
rg4 n106__vdd n108__vdd 434.8e-3
rg6 n108__vdd n110__vdd 434.8e-3
rg8 n110__vdd n112__vdd 434.8e-3
rg10 n112__vdd n114__vdd 434.8e-3
rg12 n114__vdd n116__vdd 434.8e-3
rg14 n116__vdd n118__vdd 434.8e-3
rg16 n118__vdd n120__vdd 434.8e-3
rg18 n120__vdd n122__vdd 434.8e-3
rg20 n122__vdd n105__vdd 434.8e-3
rg22 n86__vdd n106__vdd 12.5e-3
rg23 n88__vdd n108__vdd 12.5e-3
rg24 n90__vdd n110__vdd 12.5e-3
rg25 n92__vdd n112__vdd 12.5e-3
rg26 n94__vdd n114__vdd 12.5e-3
rg27 n96__vdd n116__vdd 12.5e-3
rg28 n98__vdd n118__vdd 12.5e-3
rg29 n100__vdd n120__vdd 12.5e-3
rg30 n102__vdd n122__vdd 12.5e-3
rg31 i5__r2 n2__i5__r2 333.3e-3
rg32 n7__clk_out clk_out 149.3e-3
rg33 n8__i5__r1 n9__i5__r1 250e-3
rg34 n14__i5__r2 n13__i5__r2 125e-3
rg35 n14__i5__r1 n15__i5__r1 166.7e-3
rg36 n64__reset n66__reset 933.9e-3
rg37 n66__reset n13__reset 7.8273
rg38 n66__reset n67__reset 553.4e-3
rg39 n17__i5__r0 n16__i5__r0 166.7e-3
rg40 n99__i5__clk4 n21__i5__clk4 14.1972
rg41 n40__i5__i8__net2 n19__i5__i8__net2 2.8107
rg43 n403__vdd n405__vdd 434.8e-3
rg45 n405__vdd n407__vdd 434.8e-3
rg47 n407__vdd n409__vdd 434.8e-3
rg49 n409__vdd n411__vdd 434.8e-3
rg50 n411__vdd n402__vdd 12.5e-3
rg51 n394__vdd n403__vdd 12.5e-3
rg52 n396__vdd n405__vdd 12.5e-3
rg53 n398__vdd n407__vdd 12.5e-3
rg54 n400__vdd n409__vdd 12.5e-3
rg56 n1781__vss n1783__vss 237.5e-3
rg58 n1783__vss n1785__vss 237.5e-3
rg60 n1785__vss n1787__vss 237.5e-3
rg62 n1787__vss n1789__vss 237.5e-3
rg64 n1789__vss n1791__vss 237.5e-3
rg66 n1791__vss n1793__vss 237.5e-3
rg68 n1793__vss n1795__vss 237.5e-3
rg70 n1795__vss n1797__vss 237.5e-3
rg72 n1797__vss n1799__vss 237.5e-3
rg74 n1799__vss n1801__vss 237.5e-3
rg76 n1801__vss n1803__vss 237.5e-3
rg78 n1803__vss n1805__vss 237.5e-3
rg80 n1805__vss n1807__vss 237.5e-3
rg82 n1807__vss n1809__vss 237.5e-3
rg84 n1809__vss n1811__vss 237.5e-3
rg86 n1811__vss n1458__vss 237.5e-3
rg87 n1458__vss n1547__vss 8.333e-3
rg88 n1781__vss n1813__vss 179.6e-3
rg90 n1813__vss n1815__vss 33.46e-3
rg91 n1815__vss n1816__vss 285.9e-3
rg92 n1816__vss n1817__vss 247.1e-3
rg93 n1471__vss n1781__vss 8.333e-3
rg94 n1425__vss n1781__vss 8.333e-3
rg95 n1427__vss n1783__vss 8.333e-3
rg96 n1477__vss n1783__vss 8.333e-3
rg97 n1479__vss n1785__vss 8.333e-3
rg98 n1429__vss n1785__vss 8.333e-3
rg99 n1485__vss n1787__vss 8.333e-3
rg100 n1431__vss n1787__vss 8.333e-3
rg101 n1433__vss n1789__vss 8.333e-3
rg102 n1491__vss n1789__vss 8.333e-3
rg103 n1435__vss n1791__vss 8.333e-3
rg104 n1497__vss n1791__vss 8.333e-3
rg105 n1437__vss n1793__vss 8.333e-3
rg106 n1499__vss n1793__vss 8.333e-3
rg107 n1439__vss n1795__vss 8.333e-3
rg108 n1505__vss n1795__vss 8.333e-3
rg109 n1441__vss n1797__vss 8.333e-3
rg110 n1511__vss n1797__vss 8.333e-3
rg111 n1443__vss n1799__vss 8.333e-3
rg112 n1514__vss n1799__vss 8.333e-3
rg113 n1445__vss n1801__vss 8.333e-3
rg114 n1519__vss n1801__vss 8.333e-3
rg115 n1525__vss n1803__vss 8.333e-3
rg116 n1447__vss n1803__vss 8.333e-3
rg117 n1449__vss n1805__vss 8.333e-3
rg118 n1531__vss n1805__vss 8.333e-3
rg119 n1451__vss n1807__vss 8.333e-3
rg120 n1534__vss n1807__vss 8.333e-3
rg121 n1539__vss n1809__vss 8.333e-3
rg122 n1453__vss n1809__vss 8.333e-3
rg123 n1545__vss n1811__vss 8.333e-3
rg124 n1455__vss n1811__vss 8.333e-3
rg125 n1423__vss n1813__vss 16.67e-3
rg126 n1461__vss n1813__vss 16.67e-3
rg127 n1459__vss n1815__vss 13.89e-3
rg128 n1818__vss n1819__vss 91.74e-3
rg129 n1819__vss n1820__vss 104.7e-3
rg131 n1819__vss n1822__vss 152.8e-3
rg132 n1820__vss n1823__vss 164.4e-3
rg133 n1823__vss n1824__vss 91.31e-3
rg135 n1824__vss n1826__vss 140.8e-3
rg136 n1826__vss n1827__vss 152.8e-3
rg137 n1822__vss n1463__vss 307e-3
rg138 n1820__vss n1828__vss 152.6e-3
rg139 n1828__vss n1465__vss 305e-3
rg140 n1820__vss n1829__vss 92.51e-3
rg141 n1823__vss n1830__vss 152.1e-3
rg142 n1823__vss n1831__vss 91.03e-3
rg143 n1826__vss n1832__vss 91.74e-3
rg144 n1827__vss n1469__vss 307e-3
rg145 n1830__vss n1467__vss 307e-3
rg146 n1773__vss n1820__vss 8.333e-3
rg147 n1775__vss n1824__vss 8.333e-3
rg149 n1833__vss n1835__vss 206.9e-3
rg151 n1835__vss n1837__vss 275.9e-3
rg152 n1837__vss n1838__vss 8.333e-3
rg153 n1776__vss n1833__vss 16.67e-3
rg154 n1778__vss n1835__vss 8.333e-3
rg155 n1780__vss n1837__vss 8.333e-3
rg156 n1983__vddio n1984__vddio 12.68e-3
rg157 n1984__vddio n1985__vddio 206.9e-3
rg158 n1985__vddio n1986__vddio 118.9e-3
rg159 n1986__vddio n1987__vddio 129.7e-3
rg160 n1987__vddio n1988__vddio 207.1e-3
rg161 n1988__vddio n1989__vddio 27.84e-3
rg162 n1989__vddio n1990__vddio 275.9e-3
rg163 n1990__vddio n1991__vddio 16.91e-3
rg164 n1991__vddio n1992__vddio 228.7e-3
rg165 n1992__vddio n1993__vddio 148.4e-3
rg166 n1993__vddio n1994__vddio 100.1e-3
rg167 n1994__vddio n1995__vddio 208e-3
rg168 n1995__vddio n1996__vddio 27.35e-3
rg169 n1996__vddio n1997__vddio 275.9e-3
rg170 n1997__vddio n1998__vddio 17.4e-3
rg171 n1998__vddio n1999__vddio 227.8e-3
rg172 n1999__vddio n2000__vddio 149.4e-3
rg173 n2000__vddio n2001__vddio 99.15e-3
rg174 n2001__vddio n2002__vddio 258.3e-3
rg175 n2002__vddio n2003__vddio 1.989e-3
rg176 n2003__vddio n2004__vddio 264.2e-3
rg177 n2004__vddio n799__vddio 71.06e-3
rg178 n799__vddio n2005__vddio 177.5e-3
rg179 n2005__vddio n2006__vddio 199.7e-3
rg180 n2006__vddio n2007__vddio 48.89e-3
rg181 n2007__vddio n2008__vddio 259.3e-3
rg182 n2008__vddio n2009__vddio 1.492e-3
rg183 n2009__vddio n2010__vddio 263.7e-3
rg184 n2010__vddio n2011__vddio 72.05e-3
rg185 n2011__vddio n2012__vddio 176.5e-3
rg186 n2012__vddio n2013__vddio 200.7e-3
rg187 n2013__vddio n2014__vddio 47.91e-3
rg188 n2014__vddio n203__vddio 262.7e-3
rg190 n203__vddio n2016__vddio 261.3e-3
rg191 n2016__vddio n67__vddio 114.4e-3
rg192 n1942__vddio n1984__vddio 16.67e-3
rg193 n1944__vddio n1985__vddio 8.333e-3
rg194 n1946__vddio n1987__vddio 8.333e-3
rg195 n1726__vddio n1988__vddio 13.89e-3
rg196 n1948__vddio n1989__vddio 8.333e-3
rg197 n1950__vddio n1990__vddio 8.333e-3
rg198 n1668__vddio n1991__vddio 13.89e-3
rg199 n1952__vddio n1992__vddio 8.333e-3
rg200 n1399__vddio n1993__vddio 13.89e-3
rg201 n1954__vddio n1994__vddio 8.333e-3
rg202 n1286__vddio n1995__vddio 13.89e-3
rg203 n1956__vddio n1996__vddio 8.333e-3
rg204 n1958__vddio n1997__vddio 8.333e-3
rg205 n1169__vddio n1998__vddio 13.89e-3
rg206 n1960__vddio n1999__vddio 8.333e-3
rg207 n1032__vddio n2000__vddio 13.89e-3
rg208 n1962__vddio n2001__vddio 8.333e-3
rg209 n904__vddio n2002__vddio 13.89e-3
rg210 n1964__vddio n2003__vddio 8.333e-3
rg211 n1966__vddio n2004__vddio 8.333e-3
rg212 n1968__vddio n2005__vddio 8.333e-3
rg213 n639__vddio n2006__vddio 13.89e-3
rg214 n1970__vddio n2007__vddio 8.333e-3
rg215 n568__vddio n2008__vddio 13.89e-3
rg216 n1972__vddio n2009__vddio 8.333e-3
rg217 n1974__vddio n2010__vddio 8.333e-3
rg218 n423__vddio n2011__vddio 13.89e-3
rg219 n1976__vddio n2012__vddio 8.333e-3
rg220 n273__vddio n2013__vddio 13.89e-3
rg221 n1978__vddio n2014__vddio 8.333e-3
rg222 n1980__vddio n203__vddio 8.333e-3
rg223 n1982__vddio n2016__vddio 8.333e-3
rh1 n20__i5__clk4 n21__i5__clk4 250e-3
rh2 reset n13__reset 390.8e-3
rh3 n13__reset n14__reset 605.7e-3
rh4 reset n15__reset 860.6e-3
rh5 n13__i5__i7__y2out n10__i5__i7__y2out 1.9265
rh6 n7__i5__i7__x1out n11__i5__i7__x1out 4.0994
rh7 n15__i5__i7__y1out n7__i5__i7__y1out 4.338
rh8 n12__i5__i7__x2out n10__i5__i7__x2out 2.4217
rh9 n7__i5__i7__y0out n14__i5__i7__y0out 7.8564
rh10 n12__i5__i7__x3out n10__i5__i7__x3out 2.1967
rh11 n11__i5__i7__x0out n7__i5__i7__x0out 6.4995
rh12 n1484__chipdriverout n1443__chipdriverout 22.12e-3
rh13 n1484__chipdriverout n1485__chipdriverout 92.39e-3
rh14 n1485__chipdriverout n1486__chipdriverout 87.85e-3
rh15 n1486__chipdriverout n1487__chipdriverout 92.39e-3
rh16 n1487__chipdriverout n1488__chipdriverout 87.85e-3
rh17 n1488__chipdriverout n1489__chipdriverout 91.64e-3
rh18 n1489__chipdriverout n1490__chipdriverout 88.61e-3
rh19 n1490__chipdriverout n1491__chipdriverout 141.3e-3
rh20 n1443__chipdriverout n1492__chipdriverout 142.9e-3
rh21 n1492__chipdriverout n1493__chipdriverout 91.26e-3
rh22 n1493__chipdriverout n1494__chipdriverout 91.26e-3
rh23 n1494__chipdriverout n1495__chipdriverout 85.96e-3
rh24 n1495__chipdriverout n1496__chipdriverout 140.9e-3
rh25 i5__r0 n2__i5__r0 616.8e-3
rh27 n86__vdd n88__vdd 434.9e-3
rh29 n88__vdd n90__vdd 434.9e-3
rh31 n90__vdd n92__vdd 434.9e-3
rh33 n92__vdd n94__vdd 434.9e-3
rh35 n94__vdd n96__vdd 434.9e-3
rh37 n96__vdd n98__vdd 434.9e-3
rh39 n98__vdd n100__vdd 434.9e-3
rh41 n100__vdd n102__vdd 434.9e-3
rh43 n102__vdd n104__vdd 434.9e-3
rh44 n104__vdd n105__vdd 12.5e-3
rh45 n67__vdd n86__vdd 12.5e-3
rh46 n69__vdd n88__vdd 12.5e-3
rh47 n71__vdd n90__vdd 12.5e-3
rh48 n73__vdd n92__vdd 12.5e-3
rh49 n75__vdd n94__vdd 12.5e-3
rh50 n77__vdd n96__vdd 12.5e-3
rh51 n79__vdd n98__vdd 12.5e-3
rh52 n81__vdd n100__vdd 12.5e-3
rh53 n83__vdd n102__vdd 12.5e-3
rh54 n66__vdd n104__vdd 12.5e-3
rh56 n7__i5__r1 n8__i5__r1 2.541
rh57 n13__i5__r2 n12__i5__r2 125e-3
rh58 n7__clk_out n10__clk_out 1.0003
rh59 n13__i5__r1 n14__i5__r1 333.3e-3
rh60 n778__i1__i14__net1 n779__i1__i14__net1 156.7e-3
rh61 n779__i1__i14__net1 n780__i1__i14__net1 114e-3
rh62 n780__i1__i14__net1 n781__i1__i14__net1 116e-3
rh63 n781__i1__i14__net1 n782__i1__i14__net1 114e-3
rh64 n782__i1__i14__net1 n777__i1__i14__net1 125.1e-3
rh65 n777__i1__i14__net1 n783__i1__i14__net1 94.14e-3
rh66 n783__i1__i14__net1 n784__i1__i14__net1 114e-3
rh67 n784__i1__i14__net1 n785__i1__i14__net1 113.1e-3
rh68 n785__i1__i14__net1 n786__i1__i14__net1 114e-3
rh69 n786__i1__i14__net1 n787__i1__i14__net1 116.9e-3
rh70 n787__i1__i14__net1 n788__i1__i14__net1 116.9e-3
rh71 n788__i1__i14__net1 n789__i1__i14__net1 110.2e-3
rh72 n789__i1__i14__net1 n790__i1__i14__net1 161.5e-3
rh73 n64__reset n55__reset 501.2e-3
rh74 n18__i5__i8__net2 n19__i5__i8__net2 250e-3
rh75 n15__i5__r0 n16__i5__r0 166.7e-3
rh76 n25__i5__i8__net1 n10__i5__i8__net1 1.8635
rh77 n43__i5__i6__net31 n46__i5__i6__net31 2.6155
rh78 n46__i5__i6__net31 n47__i5__i6__net31 2.4195
rh79 n47__i5__i6__net31 n16__i5__i6__net31 1.6371
rh80 n46__i5__i6__net31 n31__i5__i6__net31 185.2e-3
rh81 n47__i5__i6__net31 n23__i5__i6__net31 185.2e-3
rh82 n72__reset n52__reset 2.3976
rh83 n52__reset n67__reset 1.0519
rh84 n67__reset n42__reset 1.3152
rh85 n41__shift n42__shift 4.7996
rh86 n42__shift n14__shift 95.57e-3
rh87 n42__shift n43__shift 2.3714
rh88 n43__shift n27__shift 166.9e-3
rh89 n43__shift n37__shift 2.5972
rh90 n19__i5__i8__net5 n10__i5__i8__net5 1.8058
rh92 n39__i5__i8__net2 n40__i5__i8__net2 250e-3
rh94 n394__vdd n396__vdd 434.9e-3
rh96 n396__vdd n398__vdd 434.9e-3
rh98 n398__vdd n400__vdd 434.9e-3
rh100 n400__vdd n402__vdd 434.9e-3
rh101 n402__vdd n393__vdd 12.5e-3
rh102 n385__vdd n394__vdd 12.5e-3
rh103 n387__vdd n396__vdd 12.5e-3
rh104 n389__vdd n398__vdd 12.5e-3
rh105 n391__vdd n400__vdd 12.5e-3
rh107 n1423__vss n1425__vss 206.9e-3
rh109 n1425__vss n1427__vss 275.9e-3
rh111 n1427__vss n1429__vss 275.9e-3
rh113 n1429__vss n1431__vss 275.9e-3
rh115 n1431__vss n1433__vss 275.9e-3
rh117 n1433__vss n1435__vss 275.9e-3
rh119 n1435__vss n1437__vss 275.9e-3
rh121 n1437__vss n1439__vss 275.9e-3
rh123 n1439__vss n1441__vss 275.9e-3
rh125 n1441__vss n1443__vss 275.9e-3
rh127 n1443__vss n1445__vss 275.9e-3
rh129 n1445__vss n1447__vss 275.9e-3
rh131 n1447__vss n1449__vss 275.9e-3
rh133 n1449__vss n1451__vss 275.9e-3
rh135 n1451__vss n1453__vss 275.9e-3
rh137 n1453__vss n1455__vss 275.9e-3
rh139 n1455__vss n1457__vss 275.9e-3
rh140 n1457__vss n1458__vss 8.333e-3
rh141 n30__piso_out piso_out 160.2e-3
rh142 piso_out n19__piso_out 1.071
rh143 n19__piso_outinv n3__piso_outinv 1.312
rh145 n1773__vss n1775__vss 306.3e-3
rh146 n1775__vss n1753__vss 8.333e-3
rh147 n1752__vss n1773__vss 8.333e-3
rh149 n1776__vss n1778__vss 206.9e-3
rh151 n1778__vss n1780__vss 275.9e-3
rh152 n1780__vss n1713__vss 8.333e-3
rh153 n1713__vss n1776__vss 16.67e-3
rh154 n1713__vss n1778__vss 8.333e-3
rh156 n1942__vddio n1944__vddio 206.9e-3
rh158 n1944__vddio n1946__vddio 275.9e-3
rh160 n1946__vddio n1948__vddio 235.9e-3
rh162 n1948__vddio n1950__vddio 275.9e-3
rh164 n1950__vddio n1952__vddio 275.9e-3
rh166 n1952__vddio n1954__vddio 275.9e-3
rh168 n1954__vddio n1956__vddio 275.9e-3
rh170 n1956__vddio n1958__vddio 275.9e-3
rh172 n1958__vddio n1960__vddio 275.9e-3
rh174 n1960__vddio n1962__vddio 275.9e-3
rh176 n1962__vddio n1964__vddio 275.9e-3
rh178 n1964__vddio n1966__vddio 275.9e-3
rh180 n1966__vddio n1968__vddio 275.9e-3
rh182 n1968__vddio n1970__vddio 275.9e-3
rh184 n1970__vddio n1972__vddio 275.9e-3
rh186 n1972__vddio n1974__vddio 275.9e-3
rh188 n1974__vddio n1976__vddio 275.9e-3
rh190 n1976__vddio n1978__vddio 275.9e-3
rh192 n1978__vddio n1980__vddio 275.9e-3
rh194 n1980__vddio n1982__vddio 275.9e-3
rh195 n1982__vddio n1941__vddio 8.333e-3
rh196 n1948__vddio n1737__vddio 372.2e-3
rh197 n1737__vddio n1734__vddio 223.6e-3
rh198 n1887__vddio n1942__vddio 16.67e-3
rh199 n1892__vddio n1944__vddio 8.333e-3
rh200 n1898__vddio n1946__vddio 8.333e-3
rh201 n1904__vddio n1948__vddio 8.333e-3
rh202 n1909__vddio n1950__vddio 8.333e-3
rh203 n1911__vddio n1952__vddio 8.333e-3
rh204 n1913__vddio n1954__vddio 8.333e-3
rh205 n1915__vddio n1956__vddio 8.333e-3
rh206 n1917__vddio n1958__vddio 8.333e-3
rh207 n1919__vddio n1960__vddio 8.333e-3
rh208 n1921__vddio n1962__vddio 8.333e-3
rh209 n1923__vddio n1964__vddio 8.333e-3
rh210 n1925__vddio n1966__vddio 8.333e-3
rh211 n1927__vddio n1968__vddio 8.333e-3
rh212 n1929__vddio n1970__vddio 8.333e-3
rh213 n1931__vddio n1972__vddio 8.333e-3
rh214 n1933__vddio n1974__vddio 8.333e-3
rh215 n1935__vddio n1976__vddio 8.333e-3
rh216 n1937__vddio n1978__vddio 8.333e-3
rh217 n1939__vddio n1980__vddio 8.333e-3
ri1 n19__i5__clk4 n20__i5__clk4 500e-3
ri2 x0 n8__x0 1.458e-3
ri3 n9__x0 n7__x0 1.458e-3
ri4 n8__x0 n9__x0 51.99e-3
ri5 n7__y0 y0 65.47e-3
ri6 n6__i5__i7__x0out n7__i5__i7__x0out 500e-3
ri7 n7__i5__i7__y0out n6__i5__i7__y0out 500e-3
ri8 x1 n7__x1 2.431e-3
ri9 n8__x1 n5__x1 2.431e-3
ri10 n7__x1 n8__x1 36.58e-3
ri11 y1 n5__y1 36.58e-3
ri12 n6__i5__i7__x1out n7__i5__i7__x1out 521.2e-3
ri13 n6__i5__i7__y1out n7__i5__i7__y1out 500e-3
ri14 x2 n8__x2 2.917e-3
ri15 n9__x2 n7__x2 2.917e-3
ri16 n8__x2 n9__x2 50.06e-3
ri17 n7__y2 y2 44.29e-3
ri18 n9__i5__i7__x2out n10__i5__i7__x2out 500e-3
ri19 n10__i5__i7__y2out n9__i5__i7__y2out 500e-3
ri20 x3 n7__x3 3.403e-3
ri21 n8__x3 n5__x3 3.403e-3
ri22 n7__x3 n8__x3 53.91e-3
ri23 n5__y3 y3 46.21e-3
ri24 n64__i5__clk4 n65__i5__clk4 2.039
ri25 n65__i5__clk4 n66__i5__clk4 1.5235
ri26 n66__i5__clk4 n67__i5__clk4 1.539
ri27 n67__i5__clk4 n22__i5__clk4 1.4935
ri28 n58__i5__clk4 n65__i5__clk4 500e-3
ri29 n44__i5__clk4 n66__i5__clk4 500e-3
ri30 n30__i5__clk4 n67__i5__clk4 500e-3
ri31 n30__i5__i7__i0__net1 n29__i5__i7__i0__net1 2.039
ri32 n29__i5__i7__i0__net1 n24__i5__i7__i0__net1 1.5235
ri33 n24__i5__i7__i0__net1 n15__i5__i7__i0__net1 1.539
ri34 n15__i5__i7__i0__net1 n10__i5__i7__i0__net1 935.4e-3
ri35 n68__i5__clk4 n69__i5__clk4 2.039
ri36 n69__i5__clk4 n70__i5__clk4 1.5235
ri37 n70__i5__clk4 n71__i5__clk4 1.539
ri38 n71__i5__clk4 n23__i5__clk4 1.4935
ri39 n59__i5__clk4 n69__i5__clk4 500e-3
ri40 n45__i5__clk4 n70__i5__clk4 500e-3
ri41 n31__i5__clk4 n71__i5__clk4 500e-3
ri42 n30__i5__i7__i1__net1 n29__i5__i7__i1__net1 2.039
ri43 n29__i5__i7__i1__net1 n24__i5__i7__i1__net1 1.5235
ri44 n24__i5__i7__i1__net1 n15__i5__i7__i1__net1 1.539
ri45 n15__i5__i7__i1__net1 n10__i5__i7__i1__net1 935.4e-3
ri46 n33__reset n28__reset 1.5641
ri47 n28__reset n22__reset 1.5638
ri48 n22__reset n10__reset 1.5758
ri49 n10__reset n14__reset 19.61e-3
ri50 n34__reset n30__reset 1.5641
ri51 n30__reset n23__reset 1.5607
ri52 n23__reset n11__reset 1.5758
ri53 n11__reset n15__reset 23.18e-3
ri54 n9__i5__i7__x3out n10__i5__i7__x3out 521.2e-3
ri55 n12__i5__i7__x1out n11__i5__i7__x1out 500e-3
ri56 n11__i5__i7__x2out n12__i5__i7__x2out 1
ri57 n13__i5__i7__y2out n14__i5__i7__y2out 500e-3
ri58 n13__i5__i7__y1out n15__i5__i7__y1out 1
ri59 n11__i5__i7__x0out n12__i5__i7__x0out 1
ri60 n11__i5__i7__x3out n12__i5__i7__x3out 1
ri61 n13__i5__i7__y3out n11__i5__i7__y3out 1.8249
ri62 n13__i5__i7__y0out n14__i5__i7__y0out 500e-3
ri63 n10__i5__i7__xor2 n20__i5__i7__xor2 1.4378
ri64 n20__i5__i7__xor2 n17__i5__i7__xor2 73.87e-3
ri65 n20__i5__i7__xor2 n19__i5__i7__xor2 480.4e-3
ri66 n10__i5__i7__xor1 n20__i5__i7__xor1 1.4378
ri67 n20__i5__i7__xor1 n17__i5__i7__xor1 73.87e-3
ri68 n20__i5__i7__xor1 n18__i5__i7__xor1 480.4e-3
ri69 n11__i5__i7__i5__net1 n14__i5__i7__i5__net1 615.1e-3
ri70 n11__i5__i7__i4__net1 n14__i5__i7__i4__net1 615.1e-3
ri71 n8__i5__i7__net44 n5__i5__i7__net44 960.7e-3
ri72 n11__i5__i7__net47 n6__i5__i7__net47 945.4e-3
ri73 n13__i5__i7__net51 n20__i5__i7__net51 1.8226
ri74 n20__i5__i7__net51 n17__i5__i7__net51 142.8e-3
ri75 n20__i5__i7__net51 n19__i5__i7__net51 415e-3
ri76 n8__i5__i7__i6__net1 n14__i5__i7__i6__net1 615.1e-3
ri77 n9__i5__r0 i5__r0 250e-3
ri78 n6__i5__r1 n7__i5__r1 768.4e-3
ri79 n16__i5__i6__net31 n15__i5__i6__net31 250e-3
ri80 n13__shift n14__shift 500e-3
ri82 n67__vdd n69__vdd 447.8e-3
ri84 n69__vdd n71__vdd 447.8e-3
ri86 n71__vdd n73__vdd 447.8e-3
ri88 n73__vdd n75__vdd 447.8e-3
ri90 n75__vdd n77__vdd 447.8e-3
ri92 n77__vdd n79__vdd 447.8e-3
ri94 n79__vdd n81__vdd 447.8e-3
ri96 n81__vdd n83__vdd 447.8e-3
ri98 n83__vdd n66__vdd 447.8e-3
ri100 n47__vdd n67__vdd 12.5e-3
ri101 n49__vdd n69__vdd 12.5e-3
ri102 n51__vdd n71__vdd 12.5e-3
ri103 n53__vdd n73__vdd 12.5e-3
ri104 n55__vdd n75__vdd 12.5e-3
ri105 n57__vdd n77__vdd 12.5e-3
ri106 n59__vdd n79__vdd 12.5e-3
ri107 n61__vdd n81__vdd 12.5e-3
ri108 n63__vdd n83__vdd 12.5e-3
ri109 n6__i5__r2 i5__r2 166.7e-3
ri110 n22__i5__i7__net44 n18__i5__i7__net44 2.3033
ri111 n19__i5__i7__net46 n20__i5__i7__net46 2.769
ri112 n20__i5__i7__net46 n21__i5__i7__net46 1.0091
ri113 n21__i5__i7__net46 n5__i5__i7__net46 137e-3
ri114 n20__i5__i7__net46 n12__i5__i7__net46 121.5e-3
ri116 n22__i5__i6__net31 n23__i5__i6__net31 500e-3
ri117 n28__i5__i7__i7__net1 n22__i5__i7__i7__net1 2.3938
ri118 n8__i5__r2 n12__i5__r2 125e-3
ri119 n42__reset n41__reset 250e-3
ri120 n9__clk_out n10__clk_out 250e-3
ri121 n26__shift n27__shift 500e-3
ri122 n1916__chipdriverout n1877__chipdriverout 82.59e-3
ri123 n1877__chipdriverout n1813__chipdriverout 82.59e-3
ri124 n1813__chipdriverout n1799__chipdriverout 81.41e-3
ri125 n1799__chipdriverout n1760__chipdriverout 83.77e-3
ri126 n1760__chipdriverout n1721__chipdriverout 82.59e-3
ri127 n1721__chipdriverout n1682__chipdriverout 81.41e-3
ri128 n1682__chipdriverout n1643__chipdriverout 82.59e-3
ri129 n1643__chipdriverout n1604__chipdriverout 81.41e-3
ri130 n1604__chipdriverout n1564__chipdriverout 82.59e-3
ri131 n1564__chipdriverout n1524__chipdriverout 82.59e-3
ri132 n1524__chipdriverout n1445__chipdriverout 82.59e-3
ri133 n1445__chipdriverout n1496__chipdriverout 44.25e-3
ri134 n1496__chipdriverout n1430__chipdriverout 38.35e-3
ri135 n1430__chipdriverout n1391__chipdriverout 82.59e-3
ri136 n1391__chipdriverout n1352__chipdriverout 82.59e-3
ri137 n1352__chipdriverout n1313__chipdriverout 84.95e-3
ri138 n1313__chipdriverout n1274__chipdriverout 81.41e-3
ri139 n1274__chipdriverout n1235__chipdriverout 81.41e-3
ri140 n1235__chipdriverout n1196__chipdriverout 82.59e-3
ri141 n1196__chipdriverout n1157__chipdriverout 84.95e-3
ri142 n1157__chipdriverout n1092__chipdriverout 82.59e-3
ri143 n1092__chipdriverout n1079__chipdriverout 80.23e-3
ri144 n1079__chipdriverout n1040__chipdriverout 82.59e-3
ri145 n1040__chipdriverout n975__chipdriverout 84.95e-3
ri146 n975__chipdriverout n962__chipdriverout 81.41e-3
ri147 n962__chipdriverout n923__chipdriverout 83.77e-3
ri148 n923__chipdriverout n892__chipdriverout 81.41e-3
ri149 n892__chipdriverout n845__chipdriverout 82.59e-3
ri150 n845__chipdriverout n806__chipdriverout 82.59e-3
ri151 n806__chipdriverout n767__chipdriverout 82.59e-3
ri152 n767__chipdriverout n728__chipdriverout 84.95e-3
ri153 n728__chipdriverout n689__chipdriverout 81.41e-3
ri154 n689__chipdriverout n650__chipdriverout 82.59e-3
ri155 n650__chipdriverout n611__chipdriverout 82.59e-3
ri156 n611__chipdriverout n547__chipdriverout 82.59e-3
ri157 n547__chipdriverout n508__chipdriverout 82.59e-3
ri158 n508__chipdriverout n494__chipdriverout 82.59e-3
ri159 n494__chipdriverout n455__chipdriverout 83.77e-3
ri160 n455__chipdriverout n416__chipdriverout 80.23e-3
ri161 n416__chipdriverout n377__chipdriverout 82.59e-3
ri162 n377__chipdriverout n338__chipdriverout 82.59e-3
ri163 n338__chipdriverout n299__chipdriverout 82.59e-3
ri164 n299__chipdriverout n260__chipdriverout 82.59e-3
ri165 n260__chipdriverout n221__chipdriverout 82.59e-3
ri166 n221__chipdriverout n182__chipdriverout 84.95e-3
ri167 n182__chipdriverout n143__chipdriverout 80.23e-3
ri168 n143__chipdriverout n104__chipdriverout 82.59e-3
ri169 n104__chipdriverout n65__chipdriverout 82.59e-3
ri170 n65__chipdriverout n26__chipdriverout 82.41e-3
ri171 n1917__chipdriverout n1878__chipdriverout 82.59e-3
ri172 n1878__chipdriverout n1814__chipdriverout 82.59e-3
ri173 n1814__chipdriverout n1800__chipdriverout 81.41e-3
ri174 n1800__chipdriverout n1761__chipdriverout 83.77e-3
ri175 n1761__chipdriverout n1722__chipdriverout 82.59e-3
ri176 n1722__chipdriverout n1683__chipdriverout 81.41e-3
ri177 n1683__chipdriverout n1644__chipdriverout 82.59e-3
ri178 n1644__chipdriverout n1605__chipdriverout 81.41e-3
ri179 n1605__chipdriverout n1565__chipdriverout 82.59e-3
ri180 n1565__chipdriverout n1525__chipdriverout 82.59e-3
ri181 n1525__chipdriverout n1448__chipdriverout 82.59e-3
ri182 n1448__chipdriverout n1929__chipdriverout 44.25e-3
ri183 n1929__chipdriverout n1431__chipdriverout 38.35e-3
ri184 n1431__chipdriverout n1392__chipdriverout 82.59e-3
ri185 n1392__chipdriverout n1353__chipdriverout 82.59e-3
ri186 n1353__chipdriverout n1314__chipdriverout 84.95e-3
ri187 n1314__chipdriverout n1275__chipdriverout 81.41e-3
ri188 n1275__chipdriverout n1236__chipdriverout 81.41e-3
ri189 n1236__chipdriverout n1197__chipdriverout 82.59e-3
ri190 n1197__chipdriverout n1158__chipdriverout 84.95e-3
ri191 n1158__chipdriverout n1095__chipdriverout 82.59e-3
ri192 n1095__chipdriverout n1080__chipdriverout 80.23e-3
ri193 n1080__chipdriverout n1041__chipdriverout 82.59e-3
ri194 n1041__chipdriverout n978__chipdriverout 84.95e-3
ri195 n978__chipdriverout n963__chipdriverout 81.41e-3
ri196 n963__chipdriverout n924__chipdriverout 83.77e-3
ri197 n924__chipdriverout n893__chipdriverout 81.41e-3
ri198 n893__chipdriverout n846__chipdriverout 82.59e-3
ri199 n846__chipdriverout n807__chipdriverout 82.59e-3
ri200 n807__chipdriverout n768__chipdriverout 82.59e-3
ri201 n768__chipdriverout n729__chipdriverout 84.95e-3
ri202 n729__chipdriverout n690__chipdriverout 81.41e-3
ri203 n690__chipdriverout n651__chipdriverout 82.59e-3
ri204 n651__chipdriverout n612__chipdriverout 82.59e-3
ri205 n612__chipdriverout n548__chipdriverout 82.59e-3
ri206 n548__chipdriverout n509__chipdriverout 82.59e-3
ri207 n509__chipdriverout n495__chipdriverout 82.59e-3
ri208 n495__chipdriverout n456__chipdriverout 83.77e-3
ri209 n456__chipdriverout n417__chipdriverout 80.23e-3
ri210 n417__chipdriverout n378__chipdriverout 82.59e-3
ri211 n378__chipdriverout n339__chipdriverout 82.59e-3
ri212 n339__chipdriverout n300__chipdriverout 82.59e-3
ri213 n300__chipdriverout n261__chipdriverout 82.59e-3
ri214 n261__chipdriverout n222__chipdriverout 82.59e-3
ri215 n222__chipdriverout n183__chipdriverout 84.95e-3
ri216 n183__chipdriverout n144__chipdriverout 80.23e-3
ri217 n144__chipdriverout n105__chipdriverout 82.59e-3
ri218 n105__chipdriverout n66__chipdriverout 82.59e-3
ri219 n66__chipdriverout n27__chipdriverout 82.59e-3
ri220 n1495__chipdriverout n1929__chipdriverout 50e-3
ri221 n1918__chipdriverout n1879__chipdriverout 82.59e-3
ri222 n1879__chipdriverout n1817__chipdriverout 82.59e-3
ri223 n1817__chipdriverout n1801__chipdriverout 81.41e-3
ri224 n1801__chipdriverout n1762__chipdriverout 83.77e-3
ri225 n1762__chipdriverout n1723__chipdriverout 82.59e-3
ri226 n1723__chipdriverout n1684__chipdriverout 81.41e-3
ri227 n1684__chipdriverout n1645__chipdriverout 82.59e-3
ri228 n1645__chipdriverout n1606__chipdriverout 81.41e-3
ri229 n1606__chipdriverout n1566__chipdriverout 82.59e-3
ri230 n1566__chipdriverout n1526__chipdriverout 82.59e-3
ri231 n1526__chipdriverout n1449__chipdriverout 82.59e-3
ri232 n1449__chipdriverout n1930__chipdriverout 44.25e-3
ri233 n1930__chipdriverout n1432__chipdriverout 38.35e-3
ri234 n1432__chipdriverout n1393__chipdriverout 82.59e-3
ri235 n1393__chipdriverout n1354__chipdriverout 82.59e-3
ri236 n1354__chipdriverout n1315__chipdriverout 84.95e-3
ri237 n1315__chipdriverout n1276__chipdriverout 81.41e-3
ri238 n1276__chipdriverout n1237__chipdriverout 81.41e-3
ri239 n1237__chipdriverout n1198__chipdriverout 82.59e-3
ri240 n1198__chipdriverout n1159__chipdriverout 84.95e-3
ri241 n1159__chipdriverout n1096__chipdriverout 82.59e-3
ri242 n1096__chipdriverout n1081__chipdriverout 80.23e-3
ri243 n1081__chipdriverout n1042__chipdriverout 82.59e-3
ri244 n1042__chipdriverout n979__chipdriverout 84.95e-3
ri245 n979__chipdriverout n964__chipdriverout 81.41e-3
ri246 n964__chipdriverout n925__chipdriverout 83.77e-3
ri247 n925__chipdriverout n894__chipdriverout 81.41e-3
ri248 n894__chipdriverout n847__chipdriverout 82.59e-3
ri249 n847__chipdriverout n808__chipdriverout 82.59e-3
ri250 n808__chipdriverout n769__chipdriverout 82.59e-3
ri251 n769__chipdriverout n730__chipdriverout 84.95e-3
ri252 n730__chipdriverout n691__chipdriverout 81.41e-3
ri253 n691__chipdriverout n652__chipdriverout 82.59e-3
ri254 n652__chipdriverout n613__chipdriverout 82.59e-3
ri255 n613__chipdriverout n551__chipdriverout 82.59e-3
ri256 n551__chipdriverout n512__chipdriverout 82.59e-3
ri257 n512__chipdriverout n496__chipdriverout 82.59e-3
ri258 n496__chipdriverout n457__chipdriverout 83.77e-3
ri259 n457__chipdriverout n418__chipdriverout 80.23e-3
ri260 n418__chipdriverout n379__chipdriverout 82.59e-3
ri261 n379__chipdriverout n340__chipdriverout 82.59e-3
ri262 n340__chipdriverout n301__chipdriverout 82.59e-3
ri263 n301__chipdriverout n262__chipdriverout 82.59e-3
ri264 n262__chipdriverout n223__chipdriverout 82.59e-3
ri265 n223__chipdriverout n184__chipdriverout 84.95e-3
ri266 n184__chipdriverout n145__chipdriverout 80.23e-3
ri267 n145__chipdriverout n106__chipdriverout 82.59e-3
ri268 n106__chipdriverout n67__chipdriverout 82.59e-3
ri269 n67__chipdriverout n28__chipdriverout 82.59e-3
ri270 n1494__chipdriverout n1930__chipdriverout 50e-3
ri271 n1919__chipdriverout n1880__chipdriverout 82.59e-3
ri272 n1880__chipdriverout n1818__chipdriverout 82.59e-3
ri273 n1818__chipdriverout n1802__chipdriverout 81.41e-3
ri274 n1802__chipdriverout n1763__chipdriverout 83.77e-3
ri275 n1763__chipdriverout n1724__chipdriverout 82.59e-3
ri276 n1724__chipdriverout n1685__chipdriverout 81.41e-3
ri277 n1685__chipdriverout n1646__chipdriverout 82.59e-3
ri278 n1646__chipdriverout n1607__chipdriverout 81.41e-3
ri279 n1607__chipdriverout n1567__chipdriverout 82.59e-3
ri280 n1567__chipdriverout n1527__chipdriverout 82.59e-3
ri281 n1527__chipdriverout n1452__chipdriverout 82.59e-3
ri282 n1452__chipdriverout n1931__chipdriverout 44.25e-3
ri283 n1931__chipdriverout n1433__chipdriverout 38.35e-3
ri284 n1433__chipdriverout n1394__chipdriverout 82.59e-3
ri285 n1394__chipdriverout n1355__chipdriverout 82.59e-3
ri286 n1355__chipdriverout n1316__chipdriverout 84.95e-3
ri287 n1316__chipdriverout n1277__chipdriverout 81.41e-3
ri288 n1277__chipdriverout n1238__chipdriverout 81.41e-3
ri289 n1238__chipdriverout n1199__chipdriverout 82.59e-3
ri290 n1199__chipdriverout n1160__chipdriverout 84.95e-3
ri291 n1160__chipdriverout n1099__chipdriverout 82.59e-3
ri292 n1099__chipdriverout n1082__chipdriverout 80.23e-3
ri293 n1082__chipdriverout n1043__chipdriverout 82.59e-3
ri294 n1043__chipdriverout n982__chipdriverout 84.95e-3
ri295 n982__chipdriverout n965__chipdriverout 81.41e-3
ri296 n965__chipdriverout n926__chipdriverout 83.77e-3
ri297 n926__chipdriverout n895__chipdriverout 81.41e-3
ri298 n895__chipdriverout n848__chipdriverout 82.59e-3
ri299 n848__chipdriverout n809__chipdriverout 82.59e-3
ri300 n809__chipdriverout n770__chipdriverout 82.59e-3
ri301 n770__chipdriverout n731__chipdriverout 84.95e-3
ri302 n731__chipdriverout n692__chipdriverout 81.41e-3
ri303 n692__chipdriverout n653__chipdriverout 82.59e-3
ri304 n653__chipdriverout n614__chipdriverout 82.59e-3
ri305 n614__chipdriverout n552__chipdriverout 82.59e-3
ri306 n552__chipdriverout n513__chipdriverout 82.59e-3
ri307 n513__chipdriverout n497__chipdriverout 82.59e-3
ri308 n497__chipdriverout n458__chipdriverout 83.77e-3
ri309 n458__chipdriverout n419__chipdriverout 80.23e-3
ri310 n419__chipdriverout n380__chipdriverout 82.59e-3
ri311 n380__chipdriverout n341__chipdriverout 82.59e-3
ri312 n341__chipdriverout n302__chipdriverout 82.59e-3
ri313 n302__chipdriverout n263__chipdriverout 82.59e-3
ri314 n263__chipdriverout n224__chipdriverout 82.59e-3
ri315 n224__chipdriverout n185__chipdriverout 84.95e-3
ri316 n185__chipdriverout n146__chipdriverout 80.23e-3
ri317 n146__chipdriverout n107__chipdriverout 82.59e-3
ri318 n107__chipdriverout n68__chipdriverout 82.59e-3
ri319 n68__chipdriverout n29__chipdriverout 82.59e-3
ri320 n1493__chipdriverout n1931__chipdriverout 50e-3
ri321 n1920__chipdriverout n1881__chipdriverout 82.59e-3
ri322 n1881__chipdriverout n1821__chipdriverout 82.59e-3
ri323 n1821__chipdriverout n1803__chipdriverout 81.41e-3
ri324 n1803__chipdriverout n1764__chipdriverout 83.77e-3
ri325 n1764__chipdriverout n1725__chipdriverout 82.59e-3
ri326 n1725__chipdriverout n1686__chipdriverout 81.41e-3
ri327 n1686__chipdriverout n1647__chipdriverout 82.59e-3
ri328 n1647__chipdriverout n1608__chipdriverout 81.41e-3
ri329 n1608__chipdriverout n1568__chipdriverout 82.59e-3
ri330 n1568__chipdriverout n1528__chipdriverout 82.59e-3
ri331 n1528__chipdriverout n1453__chipdriverout 82.59e-3
ri332 n1453__chipdriverout n1932__chipdriverout 44.25e-3
ri333 n1932__chipdriverout n1434__chipdriverout 38.35e-3
ri334 n1434__chipdriverout n1395__chipdriverout 82.59e-3
ri335 n1395__chipdriverout n1356__chipdriverout 82.59e-3
ri336 n1356__chipdriverout n1317__chipdriverout 84.95e-3
ri337 n1317__chipdriverout n1278__chipdriverout 81.41e-3
ri338 n1278__chipdriverout n1239__chipdriverout 81.41e-3
ri339 n1239__chipdriverout n1200__chipdriverout 82.59e-3
ri340 n1200__chipdriverout n1161__chipdriverout 84.95e-3
ri341 n1161__chipdriverout n1100__chipdriverout 82.59e-3
ri342 n1100__chipdriverout n1083__chipdriverout 80.23e-3
ri343 n1083__chipdriverout n1044__chipdriverout 82.59e-3
ri344 n1044__chipdriverout n983__chipdriverout 84.95e-3
ri345 n983__chipdriverout n966__chipdriverout 81.41e-3
ri346 n966__chipdriverout n927__chipdriverout 83.77e-3
ri347 n927__chipdriverout n896__chipdriverout 81.41e-3
ri348 n896__chipdriverout n849__chipdriverout 82.59e-3
ri349 n849__chipdriverout n810__chipdriverout 82.59e-3
ri350 n810__chipdriverout n771__chipdriverout 82.59e-3
ri351 n771__chipdriverout n732__chipdriverout 84.95e-3
ri352 n732__chipdriverout n693__chipdriverout 81.41e-3
ri353 n693__chipdriverout n654__chipdriverout 82.59e-3
ri354 n654__chipdriverout n615__chipdriverout 82.59e-3
ri355 n615__chipdriverout n555__chipdriverout 82.59e-3
ri356 n555__chipdriverout n516__chipdriverout 82.59e-3
ri357 n516__chipdriverout n498__chipdriverout 82.59e-3
ri358 n498__chipdriverout n459__chipdriverout 83.77e-3
ri359 n459__chipdriverout n420__chipdriverout 80.23e-3
ri360 n420__chipdriverout n381__chipdriverout 82.59e-3
ri361 n381__chipdriverout n342__chipdriverout 82.59e-3
ri362 n342__chipdriverout n303__chipdriverout 82.59e-3
ri363 n303__chipdriverout n264__chipdriverout 82.59e-3
ri364 n264__chipdriverout n225__chipdriverout 82.59e-3
ri365 n225__chipdriverout n186__chipdriverout 84.95e-3
ri366 n186__chipdriverout n147__chipdriverout 80.23e-3
ri367 n147__chipdriverout n108__chipdriverout 82.59e-3
ri368 n108__chipdriverout n69__chipdriverout 82.59e-3
ri369 n69__chipdriverout n30__chipdriverout 82.59e-3
ri370 n1492__chipdriverout n1932__chipdriverout 50e-3
ri371 n1921__chipdriverout n1882__chipdriverout 82.59e-3
ri372 n1882__chipdriverout n1843__chipdriverout 80.23e-3
ri373 n1843__chipdriverout n1804__chipdriverout 83.77e-3
ri374 n1804__chipdriverout n1765__chipdriverout 83.77e-3
ri375 n1765__chipdriverout n1726__chipdriverout 82.59e-3
ri376 n1726__chipdriverout n1687__chipdriverout 81.41e-3
ri377 n1687__chipdriverout n1648__chipdriverout 82.59e-3
ri378 n1648__chipdriverout n1609__chipdriverout 81.41e-3
ri379 n1609__chipdriverout n1569__chipdriverout 82.59e-3
ri380 n1569__chipdriverout n1529__chipdriverout 82.59e-3
ri381 n1529__chipdriverout n1456__chipdriverout 82.59e-3
ri382 n1456__chipdriverout n1933__chipdriverout 44.25e-3
ri383 n1933__chipdriverout n1435__chipdriverout 38.35e-3
ri384 n1435__chipdriverout n1396__chipdriverout 82.59e-3
ri385 n1396__chipdriverout n1357__chipdriverout 82.59e-3
ri386 n1357__chipdriverout n1318__chipdriverout 84.95e-3
ri387 n1318__chipdriverout n1279__chipdriverout 81.41e-3
ri388 n1279__chipdriverout n1240__chipdriverout 81.41e-3
ri389 n1240__chipdriverout n1201__chipdriverout 82.59e-3
ri390 n1201__chipdriverout n1162__chipdriverout 84.95e-3
ri391 n1162__chipdriverout n1103__chipdriverout 82.59e-3
ri392 n1103__chipdriverout n1084__chipdriverout 80.23e-3
ri393 n1084__chipdriverout n1045__chipdriverout 82.59e-3
ri394 n1045__chipdriverout n986__chipdriverout 84.95e-3
ri395 n986__chipdriverout n967__chipdriverout 81.41e-3
ri396 n967__chipdriverout n928__chipdriverout 83.77e-3
ri397 n928__chipdriverout n873__chipdriverout 83.77e-3
ri398 n873__chipdriverout n850__chipdriverout 80.23e-3
ri399 n850__chipdriverout n811__chipdriverout 82.59e-3
ri400 n811__chipdriverout n772__chipdriverout 82.59e-3
ri401 n772__chipdriverout n733__chipdriverout 84.95e-3
ri402 n733__chipdriverout n694__chipdriverout 81.41e-3
ri403 n694__chipdriverout n655__chipdriverout 82.59e-3
ri404 n655__chipdriverout n616__chipdriverout 82.59e-3
ri405 n616__chipdriverout n556__chipdriverout 82.59e-3
ri406 n556__chipdriverout n517__chipdriverout 82.59e-3
ri407 n517__chipdriverout n499__chipdriverout 82.59e-3
ri408 n499__chipdriverout n460__chipdriverout 83.77e-3
ri409 n460__chipdriverout n421__chipdriverout 80.23e-3
ri410 n421__chipdriverout n382__chipdriverout 82.59e-3
ri411 n382__chipdriverout n343__chipdriverout 82.59e-3
ri412 n343__chipdriverout n304__chipdriverout 82.59e-3
ri413 n304__chipdriverout n265__chipdriverout 82.59e-3
ri414 n265__chipdriverout n226__chipdriverout 82.59e-3
ri415 n226__chipdriverout n187__chipdriverout 84.95e-3
ri416 n187__chipdriverout n148__chipdriverout 80.23e-3
ri417 n148__chipdriverout n109__chipdriverout 82.59e-3
ri418 n109__chipdriverout n70__chipdriverout 82.59e-3
ri419 n70__chipdriverout n31__chipdriverout 82.59e-3
ri420 n1484__chipdriverout n1933__chipdriverout 50e-3
ri421 n1922__chipdriverout n1883__chipdriverout 82.59e-3
ri422 n1883__chipdriverout n1844__chipdriverout 80.23e-3
ri423 n1844__chipdriverout n1805__chipdriverout 83.77e-3
ri424 n1805__chipdriverout n1766__chipdriverout 83.77e-3
ri425 n1766__chipdriverout n1727__chipdriverout 82.59e-3
ri426 n1727__chipdriverout n1688__chipdriverout 81.41e-3
ri427 n1688__chipdriverout n1649__chipdriverout 82.59e-3
ri428 n1649__chipdriverout n1610__chipdriverout 81.41e-3
ri429 n1610__chipdriverout n1570__chipdriverout 82.59e-3
ri430 n1570__chipdriverout n1530__chipdriverout 82.59e-3
ri431 n1530__chipdriverout n1457__chipdriverout 82.59e-3
ri432 n1457__chipdriverout n1934__chipdriverout 44.25e-3
ri433 n1934__chipdriverout n1436__chipdriverout 38.35e-3
ri434 n1436__chipdriverout n1397__chipdriverout 82.59e-3
ri435 n1397__chipdriverout n1358__chipdriverout 82.59e-3
ri436 n1358__chipdriverout n1319__chipdriverout 84.95e-3
ri437 n1319__chipdriverout n1280__chipdriverout 81.41e-3
ri438 n1280__chipdriverout n1241__chipdriverout 81.41e-3
ri439 n1241__chipdriverout n1202__chipdriverout 82.59e-3
ri440 n1202__chipdriverout n1163__chipdriverout 84.95e-3
ri441 n1163__chipdriverout n1104__chipdriverout 82.59e-3
ri442 n1104__chipdriverout n1085__chipdriverout 80.23e-3
ri443 n1085__chipdriverout n1046__chipdriverout 82.59e-3
ri444 n1046__chipdriverout n987__chipdriverout 84.95e-3
ri445 n987__chipdriverout n968__chipdriverout 81.41e-3
ri446 n968__chipdriverout n929__chipdriverout 83.77e-3
ri447 n929__chipdriverout n874__chipdriverout 83.77e-3
ri448 n874__chipdriverout n851__chipdriverout 80.23e-3
ri449 n851__chipdriverout n812__chipdriverout 82.59e-3
ri450 n812__chipdriverout n773__chipdriverout 82.59e-3
ri451 n773__chipdriverout n734__chipdriverout 84.95e-3
ri452 n734__chipdriverout n695__chipdriverout 81.41e-3
ri453 n695__chipdriverout n656__chipdriverout 82.59e-3
ri454 n656__chipdriverout n617__chipdriverout 82.59e-3
ri455 n617__chipdriverout n559__chipdriverout 82.59e-3
ri456 n559__chipdriverout n520__chipdriverout 82.59e-3
ri457 n520__chipdriverout n500__chipdriverout 82.59e-3
ri458 n500__chipdriverout n461__chipdriverout 83.77e-3
ri459 n461__chipdriverout n422__chipdriverout 80.23e-3
ri460 n422__chipdriverout n383__chipdriverout 82.59e-3
ri461 n383__chipdriverout n344__chipdriverout 82.59e-3
ri462 n344__chipdriverout n305__chipdriverout 82.59e-3
ri463 n305__chipdriverout n266__chipdriverout 82.59e-3
ri464 n266__chipdriverout n227__chipdriverout 82.59e-3
ri465 n227__chipdriverout n188__chipdriverout 84.95e-3
ri466 n188__chipdriverout n149__chipdriverout 80.23e-3
ri467 n149__chipdriverout n110__chipdriverout 82.59e-3
ri468 n110__chipdriverout n71__chipdriverout 82.59e-3
ri469 n71__chipdriverout n32__chipdriverout 82.59e-3
ri470 n1485__chipdriverout n1934__chipdriverout 50e-3
ri471 n1923__chipdriverout n1884__chipdriverout 82.59e-3
ri472 n1884__chipdriverout n1845__chipdriverout 80.23e-3
ri473 n1845__chipdriverout n1806__chipdriverout 83.77e-3
ri474 n1806__chipdriverout n1767__chipdriverout 83.77e-3
ri475 n1767__chipdriverout n1728__chipdriverout 82.59e-3
ri476 n1728__chipdriverout n1689__chipdriverout 81.41e-3
ri477 n1689__chipdriverout n1650__chipdriverout 82.59e-3
ri478 n1650__chipdriverout n1611__chipdriverout 81.41e-3
ri479 n1611__chipdriverout n1571__chipdriverout 82.59e-3
ri480 n1571__chipdriverout n1531__chipdriverout 82.59e-3
ri481 n1531__chipdriverout n1460__chipdriverout 82.59e-3
ri482 n1460__chipdriverout n1935__chipdriverout 44.25e-3
ri483 n1935__chipdriverout n1437__chipdriverout 38.35e-3
ri484 n1437__chipdriverout n1398__chipdriverout 82.59e-3
ri485 n1398__chipdriverout n1359__chipdriverout 82.59e-3
ri486 n1359__chipdriverout n1320__chipdriverout 84.95e-3
ri487 n1320__chipdriverout n1281__chipdriverout 81.41e-3
ri488 n1281__chipdriverout n1242__chipdriverout 81.41e-3
ri489 n1242__chipdriverout n1203__chipdriverout 82.59e-3
ri490 n1203__chipdriverout n1164__chipdriverout 84.95e-3
ri491 n1164__chipdriverout n1107__chipdriverout 82.59e-3
ri492 n1107__chipdriverout n1086__chipdriverout 80.23e-3
ri493 n1086__chipdriverout n1047__chipdriverout 82.59e-3
ri494 n1047__chipdriverout n990__chipdriverout 84.95e-3
ri495 n990__chipdriverout n969__chipdriverout 81.41e-3
ri496 n969__chipdriverout n930__chipdriverout 83.77e-3
ri497 n930__chipdriverout n875__chipdriverout 83.77e-3
ri498 n875__chipdriverout n852__chipdriverout 80.23e-3
ri499 n852__chipdriverout n813__chipdriverout 82.59e-3
ri500 n813__chipdriverout n774__chipdriverout 82.59e-3
ri501 n774__chipdriverout n735__chipdriverout 84.95e-3
ri502 n735__chipdriverout n696__chipdriverout 81.41e-3
ri503 n696__chipdriverout n657__chipdriverout 82.59e-3
ri504 n657__chipdriverout n618__chipdriverout 82.59e-3
ri505 n618__chipdriverout n560__chipdriverout 82.59e-3
ri506 n560__chipdriverout n521__chipdriverout 82.59e-3
ri507 n521__chipdriverout n501__chipdriverout 82.59e-3
ri508 n501__chipdriverout n462__chipdriverout 83.77e-3
ri509 n462__chipdriverout n423__chipdriverout 80.23e-3
ri510 n423__chipdriverout n384__chipdriverout 82.59e-3
ri511 n384__chipdriverout n345__chipdriverout 82.59e-3
ri512 n345__chipdriverout n306__chipdriverout 82.59e-3
ri513 n306__chipdriverout n267__chipdriverout 82.59e-3
ri514 n267__chipdriverout n228__chipdriverout 82.59e-3
ri515 n228__chipdriverout n189__chipdriverout 84.95e-3
ri516 n189__chipdriverout n150__chipdriverout 80.23e-3
ri517 n150__chipdriverout n111__chipdriverout 82.59e-3
ri518 n111__chipdriverout n72__chipdriverout 82.59e-3
ri519 n72__chipdriverout n33__chipdriverout 82.59e-3
ri520 n1486__chipdriverout n1935__chipdriverout 50e-3
ri521 n1924__chipdriverout n1885__chipdriverout 82.59e-3
ri522 n1885__chipdriverout n1846__chipdriverout 80.23e-3
ri523 n1846__chipdriverout n1807__chipdriverout 83.77e-3
ri524 n1807__chipdriverout n1768__chipdriverout 83.77e-3
ri525 n1768__chipdriverout n1729__chipdriverout 82.59e-3
ri526 n1729__chipdriverout n1690__chipdriverout 81.41e-3
ri527 n1690__chipdriverout n1651__chipdriverout 82.59e-3
ri528 n1651__chipdriverout n1612__chipdriverout 81.41e-3
ri529 n1612__chipdriverout n1572__chipdriverout 82.59e-3
ri530 n1572__chipdriverout n1532__chipdriverout 82.59e-3
ri531 n1532__chipdriverout n1461__chipdriverout 82.59e-3
ri532 n1461__chipdriverout n1936__chipdriverout 44.25e-3
ri533 n1936__chipdriverout n1438__chipdriverout 38.35e-3
ri534 n1438__chipdriverout n1399__chipdriverout 82.59e-3
ri535 n1399__chipdriverout n1360__chipdriverout 82.59e-3
ri536 n1360__chipdriverout n1321__chipdriverout 84.95e-3
ri537 n1321__chipdriverout n1282__chipdriverout 81.41e-3
ri538 n1282__chipdriverout n1243__chipdriverout 81.41e-3
ri539 n1243__chipdriverout n1204__chipdriverout 82.59e-3
ri540 n1204__chipdriverout n1165__chipdriverout 84.95e-3
ri541 n1165__chipdriverout n1108__chipdriverout 82.59e-3
ri542 n1108__chipdriverout n1087__chipdriverout 80.23e-3
ri543 n1087__chipdriverout n1048__chipdriverout 82.59e-3
ri544 n1048__chipdriverout n991__chipdriverout 84.95e-3
ri545 n991__chipdriverout n970__chipdriverout 81.41e-3
ri546 n970__chipdriverout n931__chipdriverout 83.77e-3
ri547 n931__chipdriverout n876__chipdriverout 83.77e-3
ri548 n876__chipdriverout n853__chipdriverout 80.23e-3
ri549 n853__chipdriverout n814__chipdriverout 82.59e-3
ri550 n814__chipdriverout n775__chipdriverout 82.59e-3
ri551 n775__chipdriverout n736__chipdriverout 84.95e-3
ri552 n736__chipdriverout n697__chipdriverout 81.41e-3
ri553 n697__chipdriverout n658__chipdriverout 82.59e-3
ri554 n658__chipdriverout n619__chipdriverout 82.59e-3
ri555 n619__chipdriverout n563__chipdriverout 82.59e-3
ri556 n563__chipdriverout n524__chipdriverout 82.59e-3
ri557 n524__chipdriverout n502__chipdriverout 82.59e-3
ri558 n502__chipdriverout n463__chipdriverout 83.77e-3
ri559 n463__chipdriverout n424__chipdriverout 80.23e-3
ri560 n424__chipdriverout n385__chipdriverout 82.59e-3
ri561 n385__chipdriverout n346__chipdriverout 82.59e-3
ri562 n346__chipdriverout n307__chipdriverout 82.59e-3
ri563 n307__chipdriverout n268__chipdriverout 82.59e-3
ri564 n268__chipdriverout n229__chipdriverout 82.59e-3
ri565 n229__chipdriverout n190__chipdriverout 84.95e-3
ri566 n190__chipdriverout n151__chipdriverout 80.23e-3
ri567 n151__chipdriverout n112__chipdriverout 82.59e-3
ri568 n112__chipdriverout n73__chipdriverout 82.59e-3
ri569 n73__chipdriverout n34__chipdriverout 82.59e-3
ri570 n1487__chipdriverout n1936__chipdriverout 50e-3
ri571 n1925__chipdriverout n1886__chipdriverout 82.59e-3
ri572 n1886__chipdriverout n1847__chipdriverout 80.23e-3
ri573 n1847__chipdriverout n1808__chipdriverout 83.77e-3
ri574 n1808__chipdriverout n1769__chipdriverout 83.77e-3
ri575 n1769__chipdriverout n1730__chipdriverout 82.59e-3
ri576 n1730__chipdriverout n1691__chipdriverout 81.41e-3
ri577 n1691__chipdriverout n1652__chipdriverout 82.59e-3
ri578 n1652__chipdriverout n1613__chipdriverout 81.41e-3
ri579 n1613__chipdriverout n1573__chipdriverout 82.59e-3
ri580 n1573__chipdriverout n1533__chipdriverout 82.59e-3
ri581 n1533__chipdriverout n1464__chipdriverout 82.59e-3
ri582 n1464__chipdriverout n1937__chipdriverout 44.25e-3
ri583 n1937__chipdriverout n1439__chipdriverout 38.35e-3
ri584 n1439__chipdriverout n1400__chipdriverout 82.59e-3
ri585 n1400__chipdriverout n1361__chipdriverout 82.59e-3
ri586 n1361__chipdriverout n1322__chipdriverout 84.95e-3
ri587 n1322__chipdriverout n1283__chipdriverout 81.41e-3
ri588 n1283__chipdriverout n1244__chipdriverout 81.41e-3
ri589 n1244__chipdriverout n1205__chipdriverout 82.59e-3
ri590 n1205__chipdriverout n1166__chipdriverout 84.95e-3
ri591 n1166__chipdriverout n1111__chipdriverout 82.59e-3
ri592 n1111__chipdriverout n1088__chipdriverout 80.23e-3
ri593 n1088__chipdriverout n1049__chipdriverout 82.59e-3
ri594 n1049__chipdriverout n994__chipdriverout 84.95e-3
ri595 n994__chipdriverout n971__chipdriverout 81.41e-3
ri596 n971__chipdriverout n932__chipdriverout 83.77e-3
ri597 n932__chipdriverout n877__chipdriverout 83.77e-3
ri598 n877__chipdriverout n854__chipdriverout 80.23e-3
ri599 n854__chipdriverout n815__chipdriverout 82.59e-3
ri600 n815__chipdriverout n776__chipdriverout 82.59e-3
ri601 n776__chipdriverout n737__chipdriverout 84.95e-3
ri602 n737__chipdriverout n698__chipdriverout 81.41e-3
ri603 n698__chipdriverout n659__chipdriverout 82.59e-3
ri604 n659__chipdriverout n620__chipdriverout 82.59e-3
ri605 n620__chipdriverout n564__chipdriverout 82.59e-3
ri606 n564__chipdriverout n525__chipdriverout 82.59e-3
ri607 n525__chipdriverout n503__chipdriverout 82.59e-3
ri608 n503__chipdriverout n464__chipdriverout 83.77e-3
ri609 n464__chipdriverout n425__chipdriverout 80.23e-3
ri610 n425__chipdriverout n386__chipdriverout 82.59e-3
ri611 n386__chipdriverout n347__chipdriverout 82.59e-3
ri612 n347__chipdriverout n308__chipdriverout 82.59e-3
ri613 n308__chipdriverout n269__chipdriverout 82.59e-3
ri614 n269__chipdriverout n230__chipdriverout 82.59e-3
ri615 n230__chipdriverout n191__chipdriverout 84.95e-3
ri616 n191__chipdriverout n152__chipdriverout 80.23e-3
ri617 n152__chipdriverout n113__chipdriverout 82.59e-3
ri618 n113__chipdriverout n74__chipdriverout 82.59e-3
ri619 n74__chipdriverout n35__chipdriverout 82.59e-3
ri620 n1488__chipdriverout n1937__chipdriverout 50e-3
ri621 n1926__chipdriverout n1887__chipdriverout 82.59e-3
ri622 n1887__chipdriverout n1848__chipdriverout 80.23e-3
ri623 n1848__chipdriverout n1809__chipdriverout 83.77e-3
ri624 n1809__chipdriverout n1770__chipdriverout 83.77e-3
ri625 n1770__chipdriverout n1731__chipdriverout 82.59e-3
ri626 n1731__chipdriverout n1692__chipdriverout 81.41e-3
ri627 n1692__chipdriverout n1653__chipdriverout 82.59e-3
ri628 n1653__chipdriverout n1614__chipdriverout 81.41e-3
ri629 n1614__chipdriverout n1574__chipdriverout 82.59e-3
ri630 n1574__chipdriverout n1534__chipdriverout 82.59e-3
ri631 n1534__chipdriverout n1465__chipdriverout 82.59e-3
ri632 n1465__chipdriverout n1938__chipdriverout 44.25e-3
ri633 n1938__chipdriverout n1440__chipdriverout 38.35e-3
ri634 n1440__chipdriverout n1401__chipdriverout 82.59e-3
ri635 n1401__chipdriverout n1362__chipdriverout 82.59e-3
ri636 n1362__chipdriverout n1323__chipdriverout 84.95e-3
ri637 n1323__chipdriverout n1284__chipdriverout 81.41e-3
ri638 n1284__chipdriverout n1245__chipdriverout 81.41e-3
ri639 n1245__chipdriverout n1206__chipdriverout 82.59e-3
ri640 n1206__chipdriverout n1167__chipdriverout 84.95e-3
ri641 n1167__chipdriverout n1112__chipdriverout 82.59e-3
ri642 n1112__chipdriverout n1089__chipdriverout 80.23e-3
ri643 n1089__chipdriverout n1050__chipdriverout 82.59e-3
ri644 n1050__chipdriverout n995__chipdriverout 84.95e-3
ri645 n995__chipdriverout n972__chipdriverout 81.41e-3
ri646 n972__chipdriverout n933__chipdriverout 83.77e-3
ri647 n933__chipdriverout n878__chipdriverout 83.77e-3
ri648 n878__chipdriverout n855__chipdriverout 80.23e-3
ri649 n855__chipdriverout n816__chipdriverout 82.59e-3
ri650 n816__chipdriverout n777__chipdriverout 82.59e-3
ri651 n777__chipdriverout n738__chipdriverout 84.95e-3
ri652 n738__chipdriverout n699__chipdriverout 81.41e-3
ri653 n699__chipdriverout n660__chipdriverout 82.59e-3
ri654 n660__chipdriverout n621__chipdriverout 82.59e-3
ri655 n621__chipdriverout n567__chipdriverout 82.59e-3
ri656 n567__chipdriverout n528__chipdriverout 82.59e-3
ri657 n528__chipdriverout n504__chipdriverout 82.59e-3
ri658 n504__chipdriverout n465__chipdriverout 83.77e-3
ri659 n465__chipdriverout n426__chipdriverout 80.23e-3
ri660 n426__chipdriverout n387__chipdriverout 82.59e-3
ri661 n387__chipdriverout n348__chipdriverout 82.59e-3
ri662 n348__chipdriverout n309__chipdriverout 82.59e-3
ri663 n309__chipdriverout n270__chipdriverout 82.59e-3
ri664 n270__chipdriverout n231__chipdriverout 82.59e-3
ri665 n231__chipdriverout n192__chipdriverout 84.95e-3
ri666 n192__chipdriverout n153__chipdriverout 80.23e-3
ri667 n153__chipdriverout n114__chipdriverout 82.59e-3
ri668 n114__chipdriverout n75__chipdriverout 82.59e-3
ri669 n75__chipdriverout n36__chipdriverout 82.59e-3
ri670 n1489__chipdriverout n1938__chipdriverout 50e-3
ri671 n1927__chipdriverout n1888__chipdriverout 82.59e-3
ri672 n1888__chipdriverout n1849__chipdriverout 80.23e-3
ri673 n1849__chipdriverout n1810__chipdriverout 83.77e-3
ri674 n1810__chipdriverout n1771__chipdriverout 83.77e-3
ri675 n1771__chipdriverout n1732__chipdriverout 82.59e-3
ri676 n1732__chipdriverout n1693__chipdriverout 81.41e-3
ri677 n1693__chipdriverout n1654__chipdriverout 82.59e-3
ri678 n1654__chipdriverout n1615__chipdriverout 81.41e-3
ri679 n1615__chipdriverout n1575__chipdriverout 82.59e-3
ri680 n1575__chipdriverout n1535__chipdriverout 82.59e-3
ri681 n1535__chipdriverout n1468__chipdriverout 82.59e-3
ri682 n1468__chipdriverout n1939__chipdriverout 44.25e-3
ri683 n1939__chipdriverout n1441__chipdriverout 38.35e-3
ri684 n1441__chipdriverout n1402__chipdriverout 82.59e-3
ri685 n1402__chipdriverout n1363__chipdriverout 82.59e-3
ri686 n1363__chipdriverout n1324__chipdriverout 84.95e-3
ri687 n1324__chipdriverout n1285__chipdriverout 81.41e-3
ri688 n1285__chipdriverout n1246__chipdriverout 81.41e-3
ri689 n1246__chipdriverout n1207__chipdriverout 82.59e-3
ri690 n1207__chipdriverout n1168__chipdriverout 84.95e-3
ri691 n1168__chipdriverout n1115__chipdriverout 82.59e-3
ri692 n1115__chipdriverout n1090__chipdriverout 80.23e-3
ri693 n1090__chipdriverout n1051__chipdriverout 82.59e-3
ri694 n1051__chipdriverout n998__chipdriverout 84.95e-3
ri695 n998__chipdriverout n973__chipdriverout 81.41e-3
ri696 n973__chipdriverout n934__chipdriverout 83.77e-3
ri697 n934__chipdriverout n879__chipdriverout 83.77e-3
ri698 n879__chipdriverout n856__chipdriverout 80.23e-3
ri699 n856__chipdriverout n817__chipdriverout 82.59e-3
ri700 n817__chipdriverout n778__chipdriverout 82.59e-3
ri701 n778__chipdriverout n739__chipdriverout 84.95e-3
ri702 n739__chipdriverout n700__chipdriverout 81.41e-3
ri703 n700__chipdriverout n661__chipdriverout 82.59e-3
ri704 n661__chipdriverout n622__chipdriverout 82.59e-3
ri705 n622__chipdriverout n568__chipdriverout 82.59e-3
ri706 n568__chipdriverout n529__chipdriverout 82.59e-3
ri707 n529__chipdriverout n505__chipdriverout 82.59e-3
ri708 n505__chipdriverout n466__chipdriverout 83.77e-3
ri709 n466__chipdriverout n427__chipdriverout 80.23e-3
ri710 n427__chipdriverout n388__chipdriverout 82.59e-3
ri711 n388__chipdriverout n349__chipdriverout 82.59e-3
ri712 n349__chipdriverout n310__chipdriverout 82.59e-3
ri713 n310__chipdriverout n271__chipdriverout 82.59e-3
ri714 n271__chipdriverout n232__chipdriverout 82.59e-3
ri715 n232__chipdriverout n193__chipdriverout 84.95e-3
ri716 n193__chipdriverout n154__chipdriverout 80.23e-3
ri717 n154__chipdriverout n115__chipdriverout 82.59e-3
ri718 n115__chipdriverout n76__chipdriverout 82.59e-3
ri719 n76__chipdriverout n37__chipdriverout 82.59e-3
ri720 n1490__chipdriverout n1939__chipdriverout 50e-3
ri721 n1928__chipdriverout n1889__chipdriverout 82.59e-3
ri722 n1889__chipdriverout n1850__chipdriverout 80.23e-3
ri723 n1850__chipdriverout n1811__chipdriverout 83.77e-3
ri724 n1811__chipdriverout n1772__chipdriverout 83.77e-3
ri725 n1772__chipdriverout n1733__chipdriverout 82.59e-3
ri726 n1733__chipdriverout n1694__chipdriverout 81.41e-3
ri727 n1694__chipdriverout n1655__chipdriverout 82.59e-3
ri728 n1655__chipdriverout n1616__chipdriverout 81.41e-3
ri729 n1616__chipdriverout n1576__chipdriverout 82.59e-3
ri730 n1576__chipdriverout n1536__chipdriverout 82.59e-3
ri731 n1536__chipdriverout n1469__chipdriverout 82.59e-3
ri732 n1469__chipdriverout n1491__chipdriverout 44.25e-3
ri733 n1491__chipdriverout n1442__chipdriverout 38.35e-3
ri734 n1442__chipdriverout n1403__chipdriverout 82.59e-3
ri735 n1403__chipdriverout n1364__chipdriverout 82.59e-3
ri736 n1364__chipdriverout n1325__chipdriverout 84.95e-3
ri737 n1325__chipdriverout n1286__chipdriverout 81.41e-3
ri738 n1286__chipdriverout n1247__chipdriverout 81.41e-3
ri739 n1247__chipdriverout n1208__chipdriverout 82.59e-3
ri740 n1208__chipdriverout n1169__chipdriverout 84.95e-3
ri741 n1169__chipdriverout n1116__chipdriverout 82.59e-3
ri742 n1116__chipdriverout n1091__chipdriverout 80.23e-3
ri743 n1091__chipdriverout n1052__chipdriverout 82.59e-3
ri744 n1052__chipdriverout n999__chipdriverout 84.95e-3
ri745 n999__chipdriverout n974__chipdriverout 81.41e-3
ri746 n974__chipdriverout n935__chipdriverout 83.77e-3
ri747 n935__chipdriverout n880__chipdriverout 83.77e-3
ri748 n880__chipdriverout n857__chipdriverout 80.23e-3
ri749 n857__chipdriverout n818__chipdriverout 82.59e-3
ri750 n818__chipdriverout n779__chipdriverout 82.59e-3
ri751 n779__chipdriverout n740__chipdriverout 84.95e-3
ri752 n740__chipdriverout n701__chipdriverout 81.41e-3
ri753 n701__chipdriverout n662__chipdriverout 82.59e-3
ri754 n662__chipdriverout n623__chipdriverout 82.59e-3
ri755 n623__chipdriverout n571__chipdriverout 82.59e-3
ri756 n571__chipdriverout n532__chipdriverout 82.59e-3
ri757 n532__chipdriverout n506__chipdriverout 82.59e-3
ri758 n506__chipdriverout n467__chipdriverout 83.77e-3
ri759 n467__chipdriverout n428__chipdriverout 80.23e-3
ri760 n428__chipdriverout n389__chipdriverout 82.59e-3
ri761 n389__chipdriverout n350__chipdriverout 82.59e-3
ri762 n350__chipdriverout n311__chipdriverout 82.59e-3
ri763 n311__chipdriverout n272__chipdriverout 82.59e-3
ri764 n272__chipdriverout n233__chipdriverout 82.59e-3
ri765 n233__chipdriverout n194__chipdriverout 84.95e-3
ri766 n194__chipdriverout n155__chipdriverout 80.23e-3
ri767 n155__chipdriverout n116__chipdriverout 82.59e-3
ri768 n116__chipdriverout n77__chipdriverout 82.59e-3
ri769 n77__chipdriverout n38__chipdriverout 82.59e-3
ri770 n644__vss n651__vss 165.9e-3
ri771 n651__vss n652__vss 82.59e-3
ri772 n652__vss n653__vss 82.59e-3
ri773 n653__vss n654__vss 82.59e-3
ri774 n654__vss n655__vss 82.59e-3
ri775 n655__vss n656__vss 82.59e-3
ri776 n656__vss n657__vss 82.59e-3
ri777 n657__vss n658__vss 80.23e-3
ri778 n658__vss n659__vss 82.59e-3
ri779 n659__vss n660__vss 82.59e-3
ri780 n660__vss n661__vss 82.59e-3
ri781 n661__vss n662__vss 82.59e-3
ri782 n662__vss n663__vss 82.59e-3
ri783 n663__vss n664__vss 82.59e-3
ri784 n664__vss n665__vss 82.59e-3
ri785 n665__vss n666__vss 82.59e-3
ri786 n666__vss n667__vss 82.59e-3
ri787 n667__vss n668__vss 82.59e-3
ri788 n668__vss n669__vss 82.59e-3
ri789 n669__vss n670__vss 82.59e-3
ri790 n670__vss n671__vss 82.59e-3
ri791 n671__vss n672__vss 82.59e-3
ri792 n672__vss n673__vss 80.23e-3
ri793 n673__vss n674__vss 82.59e-3
ri794 n674__vss n675__vss 82.59e-3
ri795 n675__vss n676__vss 82.59e-3
ri796 n676__vss n677__vss 82.59e-3
ri797 n677__vss n678__vss 82.59e-3
ri798 n678__vss n679__vss 82.59e-3
ri799 n679__vss n680__vss 88.49e-3
ri800 n680__vss n681__vss 82.59e-3
ri801 n681__vss n682__vss 82.59e-3
ri802 n682__vss n683__vss 82.59e-3
ri803 n683__vss n684__vss 82.59e-3
ri804 n684__vss n685__vss 82.59e-3
ri805 n685__vss n686__vss 82.59e-3
ri806 n686__vss n687__vss 82.59e-3
ri807 n687__vss n688__vss 80.23e-3
ri808 n688__vss n689__vss 82.59e-3
ri809 n689__vss n690__vss 82.59e-3
ri810 n690__vss n691__vss 82.59e-3
ri811 n691__vss n692__vss 82.59e-3
ri812 n692__vss n693__vss 82.59e-3
ri813 n693__vss n694__vss 82.59e-3
ri814 n694__vss n695__vss 82.59e-3
ri815 n695__vss n696__vss 82.59e-3
ri816 n696__vss n697__vss 82.59e-3
ri817 n697__vss n9__vss 165.9e-3
ri818 n646__vss n627__vss 82.59e-3
ri819 n627__vss n614__vss 80.23e-3
ri820 n614__vss n601__vss 83.77e-3
ri821 n601__vss n580__vss 83.77e-3
ri822 n580__vss n575__vss 82.59e-3
ri823 n575__vss n562__vss 81.41e-3
ri824 n562__vss n543__vss 82.59e-3
ri825 n543__vss n530__vss 81.41e-3
ri826 n530__vss n517__vss 82.59e-3
ri827 n517__vss n495__vss 82.59e-3
ri828 n495__vss n491__vss 82.59e-3
ri829 n491__vss n469__vss 82.59e-3
ri830 n469__vss n465__vss 82.59e-3
ri831 n465__vss n452__vss 82.59e-3
ri832 n452__vss n431__vss 84.95e-3
ri833 n431__vss n426__vss 81.41e-3
ri834 n426__vss n413__vss 81.41e-3
ri835 n413__vss n400__vss 82.59e-3
ri836 n400__vss n378__vss 84.95e-3
ri837 n378__vss n365__vss 82.59e-3
ri838 n365__vss n361__vss 80.23e-3
ri839 n361__vss n339__vss 82.59e-3
ri840 n339__vss n326__vss 84.95e-3
ri841 n326__vss n313__vss 81.41e-3
ri842 n313__vss n300__vss 83.77e-3
ri843 n300__vss n298__vss 79.05e-3
ri844 n298__vss n283__vss 84.95e-3
ri845 n283__vss n270__vss 82.59e-3
ri846 n270__vss n248__vss 82.59e-3
ri847 n248__vss n236__vss 84.95e-3
ri848 n236__vss n223__vss 81.41e-3
ri849 n223__vss n209__vss 82.59e-3
ri850 n209__vss n196__vss 82.59e-3
ri851 n196__vss n192__vss 82.59e-3
ri852 n192__vss n170__vss 82.59e-3
ri853 n170__vss n166__vss 82.59e-3
ri854 n166__vss n153__vss 83.77e-3
ri855 n153__vss n131__vss 80.23e-3
ri856 n131__vss n127__vss 82.59e-3
ri857 n127__vss n114__vss 82.59e-3
ri858 n114__vss n101__vss 82.59e-3
ri859 n101__vss n88__vss 82.59e-3
ri860 n88__vss n75__vss 82.59e-3
ri861 n75__vss n62__vss 82.59e-3
ri862 n62__vss n49__vss 82.59e-3
ri863 n49__vss n36__vss 82.59e-3
ri864 n36__vss n23__vss 82.59e-3
ri865 n23__vss n10__vss 82.59e-3
ri866 n647__vss n628__vss 82.59e-3
ri867 n628__vss n615__vss 80.23e-3
ri868 n615__vss n602__vss 83.77e-3
ri869 n602__vss n581__vss 83.77e-3
ri870 n581__vss n576__vss 82.59e-3
ri871 n576__vss n563__vss 81.41e-3
ri872 n563__vss n544__vss 82.59e-3
ri873 n544__vss n531__vss 81.41e-3
ri874 n531__vss n518__vss 82.59e-3
ri875 n518__vss n498__vss 82.59e-3
ri876 n498__vss n492__vss 82.59e-3
ri877 n492__vss n472__vss 82.59e-3
ri878 n472__vss n466__vss 82.59e-3
ri879 n466__vss n453__vss 82.59e-3
ri880 n453__vss n432__vss 84.95e-3
ri881 n432__vss n427__vss 81.41e-3
ri882 n427__vss n414__vss 81.41e-3
ri883 n414__vss n401__vss 82.59e-3
ri884 n401__vss n381__vss 84.95e-3
ri885 n381__vss n368__vss 82.59e-3
ri886 n368__vss n362__vss 80.23e-3
ri887 n362__vss n342__vss 82.59e-3
ri888 n342__vss n329__vss 84.95e-3
ri889 n329__vss n316__vss 81.41e-3
ri890 n316__vss n303__vss 83.77e-3
ri891 n303__vss n299__vss 79.05e-3
ri892 n299__vss n284__vss 84.95e-3
ri893 n284__vss n271__vss 82.59e-3
ri894 n271__vss n251__vss 82.59e-3
ri895 n251__vss n237__vss 84.95e-3
ri896 n237__vss n224__vss 81.41e-3
ri897 n224__vss n212__vss 82.59e-3
ri898 n212__vss n199__vss 82.59e-3
ri899 n199__vss n193__vss 82.59e-3
ri900 n193__vss n173__vss 82.59e-3
ri901 n173__vss n167__vss 82.59e-3
ri902 n167__vss n154__vss 83.77e-3
ri903 n154__vss n134__vss 80.23e-3
ri904 n134__vss n128__vss 82.59e-3
ri905 n128__vss n115__vss 82.59e-3
ri906 n115__vss n102__vss 82.59e-3
ri907 n102__vss n89__vss 82.59e-3
ri908 n89__vss n76__vss 82.59e-3
ri909 n76__vss n63__vss 82.59e-3
ri910 n63__vss n50__vss 82.59e-3
ri911 n50__vss n37__vss 82.59e-3
ri912 n37__vss n24__vss 82.59e-3
ri913 n24__vss n11__vss 82.59e-3
ri914 n648__vss n629__vss 82.59e-3
ri915 n629__vss n616__vss 80.23e-3
ri916 n616__vss n603__vss 83.77e-3
ri917 n603__vss n584__vss 83.77e-3
ri918 n584__vss n577__vss 82.59e-3
ri919 n577__vss n564__vss 81.41e-3
ri920 n564__vss n545__vss 82.59e-3
ri921 n545__vss n532__vss 81.41e-3
ri922 n532__vss n519__vss 82.59e-3
ri923 n519__vss n499__vss 82.59e-3
ri924 n499__vss n493__vss 82.59e-3
ri925 n493__vss n473__vss 82.59e-3
ri926 n473__vss n467__vss 82.59e-3
ri927 n467__vss n454__vss 82.59e-3
ri928 n454__vss n435__vss 84.95e-3
ri929 n435__vss n428__vss 81.41e-3
ri930 n428__vss n415__vss 81.41e-3
ri931 n415__vss n402__vss 82.59e-3
ri932 n402__vss n382__vss 84.95e-3
ri933 n382__vss n369__vss 82.59e-3
ri934 n369__vss n363__vss 80.23e-3
ri935 n363__vss n343__vss 82.59e-3
ri936 n343__vss n330__vss 84.95e-3
ri937 n330__vss n317__vss 81.41e-3
ri938 n317__vss n304__vss 83.77e-3
ri939 n304__vss n287__vss 80.23e-3
ri940 n287__vss n285__vss 83.77e-3
ri941 n285__vss n272__vss 82.59e-3
ri942 n272__vss n252__vss 82.59e-3
ri943 n252__vss n240__vss 84.95e-3
ri944 n240__vss n227__vss 81.41e-3
ri945 n227__vss n213__vss 82.59e-3
ri946 n213__vss n200__vss 82.59e-3
ri947 n200__vss n194__vss 82.59e-3
ri948 n194__vss n174__vss 82.59e-3
ri949 n174__vss n168__vss 82.59e-3
ri950 n168__vss n155__vss 83.77e-3
ri951 n155__vss n135__vss 80.23e-3
ri952 n135__vss n129__vss 82.59e-3
ri953 n129__vss n116__vss 82.59e-3
ri954 n116__vss n103__vss 82.59e-3
ri955 n103__vss n90__vss 82.59e-3
ri956 n90__vss n77__vss 82.59e-3
ri957 n77__vss n64__vss 82.59e-3
ri958 n64__vss n51__vss 82.59e-3
ri959 n51__vss n38__vss 82.59e-3
ri960 n38__vss n25__vss 82.59e-3
ri961 n25__vss n12__vss 82.59e-3
ri962 n649__vss n630__vss 82.59e-3
ri963 n630__vss n617__vss 80.23e-3
ri964 n617__vss n604__vss 83.77e-3
ri965 n604__vss n585__vss 83.77e-3
ri966 n585__vss n578__vss 82.59e-3
ri967 n578__vss n565__vss 81.41e-3
ri968 n565__vss n546__vss 82.59e-3
ri969 n546__vss n533__vss 81.41e-3
ri970 n533__vss n520__vss 82.59e-3
ri971 n520__vss n502__vss 82.59e-3
ri972 n502__vss n494__vss 82.59e-3
ri973 n494__vss n476__vss 82.59e-3
ri974 n476__vss n468__vss 82.59e-3
ri975 n468__vss n455__vss 82.59e-3
ri976 n455__vss n436__vss 84.95e-3
ri977 n436__vss n429__vss 81.41e-3
ri978 n429__vss n416__vss 81.41e-3
ri979 n416__vss n403__vss 82.59e-3
ri980 n403__vss n385__vss 84.95e-3
ri981 n385__vss n372__vss 82.59e-3
ri982 n372__vss n364__vss 80.23e-3
ri983 n364__vss n346__vss 82.59e-3
ri984 n346__vss n333__vss 84.95e-3
ri985 n333__vss n320__vss 81.41e-3
ri986 n320__vss n307__vss 83.77e-3
ri987 n307__vss n290__vss 80.23e-3
ri988 n290__vss n286__vss 83.77e-3
ri989 n286__vss n273__vss 82.59e-3
ri990 n273__vss n255__vss 82.59e-3
ri991 n255__vss n241__vss 84.95e-3
ri992 n241__vss n228__vss 81.41e-3
ri993 n228__vss n216__vss 82.59e-3
ri994 n216__vss n203__vss 82.59e-3
ri995 n203__vss n195__vss 82.59e-3
ri996 n195__vss n177__vss 82.59e-3
ri997 n177__vss n169__vss 82.59e-3
ri998 n169__vss n156__vss 83.77e-3
ri999 n156__vss n138__vss 80.23e-3
ri1000 n138__vss n130__vss 82.59e-3
ri1001 n130__vss n117__vss 82.59e-3
ri1002 n117__vss n104__vss 82.59e-3
ri1003 n104__vss n91__vss 82.59e-3
ri1004 n91__vss n78__vss 82.59e-3
ri1005 n78__vss n65__vss 82.59e-3
ri1006 n65__vss n52__vss 82.59e-3
ri1007 n52__vss n39__vss 82.59e-3
ri1008 n39__vss n26__vss 82.59e-3
ri1009 n26__vss n13__vss 82.59e-3
ri1010 n1113__vddio n1092__vddio 82.59e-3
ri1011 n1092__vddio n1071__vddio 80.23e-3
ri1012 n1071__vddio n1050__vddio 83.77e-3
ri1013 n1050__vddio n1006__vddio 83.77e-3
ri1014 n1006__vddio n998__vddio 82.59e-3
ri1015 n998__vddio n977__vddio 81.41e-3
ri1016 n977__vddio n956__vddio 82.59e-3
ri1017 n956__vddio n935__vddio 81.41e-3
ri1018 n935__vddio n914__vddio 82.59e-3
ri1019 n914__vddio n869__vddio 82.59e-3
ri1020 n869__vddio n862__vddio 82.59e-3
ri1021 n862__vddio n827__vddio 82.59e-3
ri1022 n827__vddio n814__vddio 82.59e-3
ri1023 n814__vddio n789__vddio 82.59e-3
ri1024 n789__vddio n768__vddio 84.95e-3
ri1025 n768__vddio n747__vddio 81.41e-3
ri1026 n747__vddio n726__vddio 81.41e-3
ri1027 n726__vddio n705__vddio 82.59e-3
ri1028 n705__vddio n670__vddio 84.95e-3
ri1029 n670__vddio n663__vddio 82.59e-3
ri1030 n663__vddio n632__vddio 80.23e-3
ri1031 n632__vddio n597__vddio 82.59e-3
ri1032 n597__vddio n590__vddio 84.95e-3
ri1033 n590__vddio n545__vddio 81.41e-3
ri1034 n545__vddio n538__vddio 83.77e-3
ri1035 n538__vddio n517__vddio 83.77e-3
ri1036 n517__vddio n496__vddio 80.23e-3
ri1037 n496__vddio n475__vddio 82.59e-3
ri1038 n475__vddio n434__vddio 82.59e-3
ri1039 n434__vddio n410__vddio 84.95e-3
ri1040 n410__vddio n389__vddio 81.41e-3
ri1041 n389__vddio n367__vddio 82.59e-3
ri1042 n367__vddio n346__vddio 82.59e-3
ri1043 n346__vddio n339__vddio 82.59e-3
ri1044 n339__vddio n304__vddio 82.59e-3
ri1045 n304__vddio n297__vddio 82.59e-3
ri1046 n297__vddio n266__vddio 83.77e-3
ri1047 n266__vddio n231__vddio 80.23e-3
ri1048 n231__vddio n224__vddio 82.59e-3
ri1049 n224__vddio n193__vddio 82.59e-3
ri1050 n193__vddio n172__vddio 82.59e-3
ri1051 n172__vddio n151__vddio 82.59e-3
ri1052 n151__vddio n130__vddio 82.59e-3
ri1053 n130__vddio n109__vddio 82.59e-3
ri1054 n109__vddio n82__vddio 82.59e-3
ri1055 n82__vddio n57__vddio 82.59e-3
ri1056 n57__vddio n36__vddio 82.59e-3
ri1057 n36__vddio n15__vddio 82.59e-3
ri1058 n1114__vddio n1093__vddio 82.59e-3
ri1059 n1093__vddio n1072__vddio 80.23e-3
ri1060 n1072__vddio n1051__vddio 83.77e-3
ri1061 n1051__vddio n1007__vddio 83.77e-3
ri1062 n1007__vddio n999__vddio 82.59e-3
ri1063 n999__vddio n978__vddio 81.41e-3
ri1064 n978__vddio n957__vddio 82.59e-3
ri1065 n957__vddio n936__vddio 81.41e-3
ri1066 n936__vddio n915__vddio 82.59e-3
ri1067 n915__vddio n872__vddio 82.59e-3
ri1068 n872__vddio n863__vddio 82.59e-3
ri1069 n863__vddio n830__vddio 82.59e-3
ri1070 n830__vddio n815__vddio 82.59e-3
ri1071 n815__vddio n790__vddio 82.59e-3
ri1072 n790__vddio n769__vddio 84.95e-3
ri1073 n769__vddio n748__vddio 81.41e-3
ri1074 n748__vddio n727__vddio 81.41e-3
ri1075 n727__vddio n706__vddio 82.59e-3
ri1076 n706__vddio n673__vddio 84.95e-3
ri1077 n673__vddio n664__vddio 82.59e-3
ri1078 n664__vddio n633__vddio 80.23e-3
ri1079 n633__vddio n600__vddio 82.59e-3
ri1080 n600__vddio n591__vddio 84.95e-3
ri1081 n591__vddio n548__vddio 81.41e-3
ri1082 n548__vddio n539__vddio 83.77e-3
ri1083 n539__vddio n518__vddio 83.77e-3
ri1084 n518__vddio n497__vddio 80.23e-3
ri1085 n497__vddio n476__vddio 82.59e-3
ri1086 n476__vddio n437__vddio 82.59e-3
ri1087 n437__vddio n411__vddio 84.95e-3
ri1088 n411__vddio n390__vddio 81.41e-3
ri1089 n390__vddio n370__vddio 82.59e-3
ri1090 n370__vddio n349__vddio 82.59e-3
ri1091 n349__vddio n340__vddio 82.59e-3
ri1092 n340__vddio n307__vddio 82.59e-3
ri1093 n307__vddio n298__vddio 82.59e-3
ri1094 n298__vddio n267__vddio 83.77e-3
ri1095 n267__vddio n234__vddio 80.23e-3
ri1096 n234__vddio n225__vddio 82.59e-3
ri1097 n225__vddio n194__vddio 82.59e-3
ri1098 n194__vddio n173__vddio 82.59e-3
ri1099 n173__vddio n152__vddio 82.59e-3
ri1100 n152__vddio n131__vddio 82.59e-3
ri1101 n131__vddio n110__vddio 82.59e-3
ri1102 n110__vddio n83__vddio 82.59e-3
ri1103 n83__vddio n58__vddio 82.59e-3
ri1104 n58__vddio n37__vddio 82.59e-3
ri1105 n37__vddio n16__vddio 82.59e-3
ri1106 n1115__vddio n1094__vddio 82.59e-3
ri1107 n1094__vddio n1073__vddio 80.23e-3
ri1108 n1073__vddio n1052__vddio 83.77e-3
ri1109 n1052__vddio n1010__vddio 83.77e-3
ri1110 n1010__vddio n1000__vddio 82.59e-3
ri1111 n1000__vddio n979__vddio 81.41e-3
ri1112 n979__vddio n958__vddio 82.59e-3
ri1113 n958__vddio n937__vddio 81.41e-3
ri1114 n937__vddio n916__vddio 82.59e-3
ri1115 n916__vddio n873__vddio 82.59e-3
ri1116 n873__vddio n864__vddio 82.59e-3
ri1117 n864__vddio n831__vddio 82.59e-3
ri1118 n831__vddio n816__vddio 82.59e-3
ri1119 n816__vddio n791__vddio 82.59e-3
ri1120 n791__vddio n770__vddio 84.95e-3
ri1121 n770__vddio n749__vddio 81.41e-3
ri1122 n749__vddio n728__vddio 81.41e-3
ri1123 n728__vddio n707__vddio 82.59e-3
ri1124 n707__vddio n674__vddio 84.95e-3
ri1125 n674__vddio n665__vddio 82.59e-3
ri1126 n665__vddio n634__vddio 80.23e-3
ri1127 n634__vddio n601__vddio 82.59e-3
ri1128 n601__vddio n592__vddio 84.95e-3
ri1129 n592__vddio n549__vddio 81.41e-3
ri1130 n549__vddio n540__vddio 83.77e-3
ri1131 n540__vddio n519__vddio 83.77e-3
ri1132 n519__vddio n498__vddio 80.23e-3
ri1133 n498__vddio n477__vddio 82.59e-3
ri1134 n477__vddio n438__vddio 82.59e-3
ri1135 n438__vddio n414__vddio 84.95e-3
ri1136 n414__vddio n393__vddio 81.41e-3
ri1137 n393__vddio n371__vddio 82.59e-3
ri1138 n371__vddio n350__vddio 82.59e-3
ri1139 n350__vddio n341__vddio 82.59e-3
ri1140 n341__vddio n308__vddio 82.59e-3
ri1141 n308__vddio n299__vddio 82.59e-3
ri1142 n299__vddio n268__vddio 83.77e-3
ri1143 n268__vddio n235__vddio 80.23e-3
ri1144 n235__vddio n226__vddio 82.59e-3
ri1145 n226__vddio n195__vddio 82.59e-3
ri1146 n195__vddio n174__vddio 82.59e-3
ri1147 n174__vddio n153__vddio 82.59e-3
ri1148 n153__vddio n132__vddio 82.59e-3
ri1149 n132__vddio n111__vddio 82.59e-3
ri1150 n111__vddio n84__vddio 82.59e-3
ri1151 n84__vddio n59__vddio 82.59e-3
ri1152 n59__vddio n38__vddio 82.59e-3
ri1153 n38__vddio n17__vddio 82.59e-3
ri1154 n1116__vddio n1095__vddio 82.59e-3
ri1155 n1095__vddio n1074__vddio 80.23e-3
ri1156 n1074__vddio n1053__vddio 83.77e-3
ri1157 n1053__vddio n1011__vddio 83.77e-3
ri1158 n1011__vddio n1001__vddio 82.59e-3
ri1159 n1001__vddio n980__vddio 81.41e-3
ri1160 n980__vddio n959__vddio 82.59e-3
ri1161 n959__vddio n938__vddio 81.41e-3
ri1162 n938__vddio n917__vddio 82.59e-3
ri1163 n917__vddio n876__vddio 82.59e-3
ri1164 n876__vddio n865__vddio 82.59e-3
ri1165 n865__vddio n834__vddio 82.59e-3
ri1166 n834__vddio n817__vddio 82.59e-3
ri1167 n817__vddio n792__vddio 82.59e-3
ri1168 n792__vddio n771__vddio 84.95e-3
ri1169 n771__vddio n750__vddio 81.41e-3
ri1170 n750__vddio n729__vddio 81.41e-3
ri1171 n729__vddio n708__vddio 82.59e-3
ri1172 n708__vddio n677__vddio 84.95e-3
ri1173 n677__vddio n666__vddio 82.59e-3
ri1174 n666__vddio n635__vddio 80.23e-3
ri1175 n635__vddio n604__vddio 82.59e-3
ri1176 n604__vddio n593__vddio 84.95e-3
ri1177 n593__vddio n552__vddio 81.41e-3
ri1178 n552__vddio n541__vddio 83.77e-3
ri1179 n541__vddio n520__vddio 83.77e-3
ri1180 n520__vddio n499__vddio 80.23e-3
ri1181 n499__vddio n478__vddio 82.59e-3
ri1182 n478__vddio n441__vddio 82.59e-3
ri1183 n441__vddio n415__vddio 84.95e-3
ri1184 n415__vddio n394__vddio 81.41e-3
ri1185 n394__vddio n374__vddio 82.59e-3
ri1186 n374__vddio n353__vddio 82.59e-3
ri1187 n353__vddio n342__vddio 82.59e-3
ri1188 n342__vddio n311__vddio 82.59e-3
ri1189 n311__vddio n300__vddio 82.59e-3
ri1190 n300__vddio n269__vddio 83.77e-3
ri1191 n269__vddio n238__vddio 80.23e-3
ri1192 n238__vddio n227__vddio 82.59e-3
ri1193 n227__vddio n196__vddio 82.59e-3
ri1194 n196__vddio n175__vddio 82.59e-3
ri1195 n175__vddio n154__vddio 82.59e-3
ri1196 n154__vddio n133__vddio 82.59e-3
ri1197 n133__vddio n112__vddio 82.59e-3
ri1198 n112__vddio n85__vddio 82.59e-3
ri1199 n85__vddio n60__vddio 82.59e-3
ri1200 n60__vddio n39__vddio 82.59e-3
ri1201 n39__vddio n18__vddio 82.59e-3
ri1202 n1117__vddio n1096__vddio 82.59e-3
ri1203 n1096__vddio n1075__vddio 80.23e-3
ri1204 n1075__vddio n1054__vddio 83.77e-3
ri1205 n1054__vddio n1014__vddio 83.77e-3
ri1206 n1014__vddio n1002__vddio 82.59e-3
ri1207 n1002__vddio n981__vddio 81.41e-3
ri1208 n981__vddio n960__vddio 82.59e-3
ri1209 n960__vddio n939__vddio 81.41e-3
ri1210 n939__vddio n918__vddio 82.59e-3
ri1211 n918__vddio n877__vddio 82.59e-3
ri1212 n877__vddio n866__vddio 82.59e-3
ri1213 n866__vddio n835__vddio 82.59e-3
ri1214 n835__vddio n818__vddio 82.59e-3
ri1215 n818__vddio n793__vddio 82.59e-3
ri1216 n793__vddio n772__vddio 84.95e-3
ri1217 n772__vddio n751__vddio 81.41e-3
ri1218 n751__vddio n730__vddio 81.41e-3
ri1219 n730__vddio n709__vddio 82.59e-3
ri1220 n709__vddio n678__vddio 84.95e-3
ri1221 n678__vddio n667__vddio 82.59e-3
ri1222 n667__vddio n636__vddio 80.23e-3
ri1223 n636__vddio n605__vddio 82.59e-3
ri1224 n605__vddio n594__vddio 84.95e-3
ri1225 n594__vddio n553__vddio 81.41e-3
ri1226 n553__vddio n542__vddio 83.77e-3
ri1227 n542__vddio n521__vddio 83.77e-3
ri1228 n521__vddio n500__vddio 80.23e-3
ri1229 n500__vddio n479__vddio 82.59e-3
ri1230 n479__vddio n442__vddio 82.59e-3
ri1231 n442__vddio n418__vddio 84.95e-3
ri1232 n418__vddio n397__vddio 81.41e-3
ri1233 n397__vddio n375__vddio 82.59e-3
ri1234 n375__vddio n354__vddio 82.59e-3
ri1235 n354__vddio n343__vddio 82.59e-3
ri1236 n343__vddio n312__vddio 82.59e-3
ri1237 n312__vddio n301__vddio 82.59e-3
ri1238 n301__vddio n270__vddio 83.77e-3
ri1239 n270__vddio n239__vddio 80.23e-3
ri1240 n239__vddio n228__vddio 82.59e-3
ri1241 n228__vddio n197__vddio 82.59e-3
ri1242 n197__vddio n176__vddio 82.59e-3
ri1243 n176__vddio n155__vddio 82.59e-3
ri1244 n155__vddio n134__vddio 82.59e-3
ri1245 n134__vddio n113__vddio 82.59e-3
ri1246 n113__vddio n86__vddio 82.59e-3
ri1247 n86__vddio n61__vddio 82.59e-3
ri1248 n61__vddio n40__vddio 82.59e-3
ri1249 n40__vddio n19__vddio 82.59e-3
ri1250 n1118__vddio n1097__vddio 82.59e-3
ri1251 n1097__vddio n1076__vddio 80.23e-3
ri1252 n1076__vddio n1055__vddio 83.77e-3
ri1253 n1055__vddio n1015__vddio 83.77e-3
ri1254 n1015__vddio n1003__vddio 82.59e-3
ri1255 n1003__vddio n982__vddio 81.41e-3
ri1256 n982__vddio n961__vddio 82.59e-3
ri1257 n961__vddio n940__vddio 81.41e-3
ri1258 n940__vddio n919__vddio 82.59e-3
ri1259 n919__vddio n880__vddio 82.59e-3
ri1260 n880__vddio n867__vddio 82.59e-3
ri1261 n867__vddio n838__vddio 82.59e-3
ri1262 n838__vddio n819__vddio 82.59e-3
ri1263 n819__vddio n794__vddio 82.59e-3
ri1264 n794__vddio n773__vddio 84.95e-3
ri1265 n773__vddio n752__vddio 81.41e-3
ri1266 n752__vddio n731__vddio 81.41e-3
ri1267 n731__vddio n710__vddio 82.59e-3
ri1268 n710__vddio n681__vddio 84.95e-3
ri1269 n681__vddio n668__vddio 82.59e-3
ri1270 n668__vddio n637__vddio 80.23e-3
ri1271 n637__vddio n608__vddio 82.59e-3
ri1272 n608__vddio n595__vddio 84.95e-3
ri1273 n595__vddio n556__vddio 81.41e-3
ri1274 n556__vddio n543__vddio 83.77e-3
ri1275 n543__vddio n522__vddio 83.77e-3
ri1276 n522__vddio n501__vddio 80.23e-3
ri1277 n501__vddio n480__vddio 82.59e-3
ri1278 n480__vddio n445__vddio 82.59e-3
ri1279 n445__vddio n419__vddio 84.95e-3
ri1280 n419__vddio n398__vddio 81.41e-3
ri1281 n398__vddio n378__vddio 82.59e-3
ri1282 n378__vddio n357__vddio 82.59e-3
ri1283 n357__vddio n344__vddio 82.59e-3
ri1284 n344__vddio n315__vddio 82.59e-3
ri1285 n315__vddio n302__vddio 82.59e-3
ri1286 n302__vddio n271__vddio 83.77e-3
ri1287 n271__vddio n242__vddio 80.23e-3
ri1288 n242__vddio n229__vddio 82.59e-3
ri1289 n229__vddio n198__vddio 82.59e-3
ri1290 n198__vddio n177__vddio 82.59e-3
ri1291 n177__vddio n156__vddio 82.59e-3
ri1292 n156__vddio n135__vddio 82.59e-3
ri1293 n135__vddio n114__vddio 82.59e-3
ri1294 n114__vddio n87__vddio 82.59e-3
ri1295 n87__vddio n62__vddio 82.59e-3
ri1296 n62__vddio n41__vddio 82.59e-3
ri1297 n41__vddio n20__vddio 82.59e-3
ri1298 n1119__vddio n1098__vddio 82.59e-3
ri1299 n1098__vddio n1077__vddio 80.23e-3
ri1300 n1077__vddio n1056__vddio 83.77e-3
ri1301 n1056__vddio n1018__vddio 83.77e-3
ri1302 n1018__vddio n1004__vddio 82.59e-3
ri1303 n1004__vddio n983__vddio 81.41e-3
ri1304 n983__vddio n962__vddio 82.59e-3
ri1305 n962__vddio n941__vddio 81.41e-3
ri1306 n941__vddio n920__vddio 82.59e-3
ri1307 n920__vddio n881__vddio 82.59e-3
ri1308 n881__vddio n868__vddio 82.59e-3
ri1309 n868__vddio n839__vddio 82.59e-3
ri1310 n839__vddio n820__vddio 82.59e-3
ri1311 n820__vddio n795__vddio 82.59e-3
ri1312 n795__vddio n774__vddio 84.95e-3
ri1313 n774__vddio n753__vddio 81.41e-3
ri1314 n753__vddio n732__vddio 81.41e-3
ri1315 n732__vddio n711__vddio 82.59e-3
ri1316 n711__vddio n682__vddio 84.95e-3
ri1317 n682__vddio n669__vddio 82.59e-3
ri1318 n669__vddio n638__vddio 80.23e-3
ri1319 n638__vddio n609__vddio 82.59e-3
ri1320 n609__vddio n596__vddio 84.95e-3
ri1321 n596__vddio n557__vddio 81.41e-3
ri1322 n557__vddio n544__vddio 83.77e-3
ri1323 n544__vddio n523__vddio 83.77e-3
ri1324 n523__vddio n502__vddio 80.23e-3
ri1325 n502__vddio n481__vddio 82.59e-3
ri1326 n481__vddio n446__vddio 82.59e-3
ri1327 n446__vddio n422__vddio 84.95e-3
ri1328 n422__vddio n401__vddio 81.41e-3
ri1329 n401__vddio n379__vddio 82.59e-3
ri1330 n379__vddio n358__vddio 82.59e-3
ri1331 n358__vddio n345__vddio 82.59e-3
ri1332 n345__vddio n316__vddio 82.59e-3
ri1333 n316__vddio n303__vddio 82.59e-3
ri1334 n303__vddio n272__vddio 83.77e-3
ri1335 n272__vddio n243__vddio 80.23e-3
ri1336 n243__vddio n230__vddio 82.59e-3
ri1337 n230__vddio n199__vddio 82.59e-3
ri1338 n199__vddio n178__vddio 82.59e-3
ri1339 n178__vddio n157__vddio 82.59e-3
ri1340 n157__vddio n136__vddio 82.59e-3
ri1341 n136__vddio n115__vddio 82.59e-3
ri1342 n115__vddio n88__vddio 82.59e-3
ri1343 n88__vddio n63__vddio 82.59e-3
ri1344 n63__vddio n42__vddio 82.59e-3
ri1345 n42__vddio n21__vddio 82.59e-3
ri1346 n1112__vddio n1121__vddio 165.9e-3
ri1347 n1121__vddio n1122__vddio 80.23e-3
ri1348 n1122__vddio n1123__vddio 83.77e-3
ri1349 n1123__vddio n1124__vddio 83.77e-3
ri1350 n1124__vddio n1125__vddio 82.59e-3
ri1351 n1125__vddio n1126__vddio 81.41e-3
ri1352 n1126__vddio n1127__vddio 82.59e-3
ri1353 n1127__vddio n1128__vddio 81.41e-3
ri1354 n1128__vddio n1129__vddio 82.59e-3
ri1355 n1129__vddio n1130__vddio 82.59e-3
ri1356 n1130__vddio n1131__vddio 82.59e-3
ri1357 n1131__vddio n1132__vddio 82.59e-3
ri1358 n1132__vddio n1133__vddio 82.59e-3
ri1359 n1133__vddio n1134__vddio 82.59e-3
ri1360 n1134__vddio n1135__vddio 84.95e-3
ri1361 n1135__vddio n1136__vddio 81.41e-3
ri1362 n1136__vddio n1137__vddio 81.41e-3
ri1363 n1137__vddio n1138__vddio 82.59e-3
ri1364 n1138__vddio n1139__vddio 84.95e-3
ri1365 n1139__vddio n1140__vddio 82.59e-3
ri1366 n1140__vddio n1141__vddio 80.23e-3
ri1367 n1141__vddio n1142__vddio 82.59e-3
ri1368 n1142__vddio n1143__vddio 84.95e-3
ri1369 n1143__vddio n1144__vddio 81.41e-3
ri1370 n1144__vddio n1145__vddio 83.77e-3
ri1371 n1145__vddio n1146__vddio 83.77e-3
ri1372 n1146__vddio n1147__vddio 80.23e-3
ri1373 n1147__vddio n1148__vddio 82.59e-3
ri1374 n1148__vddio n1149__vddio 82.59e-3
ri1375 n1149__vddio n1150__vddio 84.95e-3
ri1376 n1150__vddio n1151__vddio 81.41e-3
ri1377 n1151__vddio n1152__vddio 82.59e-3
ri1378 n1152__vddio n1153__vddio 82.59e-3
ri1379 n1153__vddio n1154__vddio 82.59e-3
ri1380 n1154__vddio n1155__vddio 82.59e-3
ri1381 n1155__vddio n1156__vddio 82.59e-3
ri1382 n1156__vddio n1157__vddio 83.77e-3
ri1383 n1157__vddio n1158__vddio 80.23e-3
ri1384 n1158__vddio n1159__vddio 82.59e-3
ri1385 n1159__vddio n1160__vddio 82.59e-3
ri1386 n1160__vddio n1161__vddio 82.59e-3
ri1387 n1161__vddio n1162__vddio 82.59e-3
ri1388 n1162__vddio n1163__vddio 82.59e-3
ri1389 n1163__vddio n1164__vddio 82.59e-3
ri1390 n1164__vddio n1165__vddio 82.59e-3
ri1391 n1165__vddio n1166__vddio 82.59e-3
ri1392 n1166__vddio n1167__vddio 82.59e-3
ri1393 n1167__vddio n14__vddio 165.9e-3
ri1394 n13__i5__r1 n16__i5__r1 166.7e-3
ri1395 n777__i1__i14__net1 n775__i1__i14__net1 130.2e-3
ri1397 n775__i1__i14__net1 n771__i1__i14__net1 18.86e-3
ri1399 n771__i1__i14__net1 n767__i1__i14__net1 22.45e-3
ri1401 n767__i1__i14__net1 n762__i1__i14__net1 18.86e-3
ri1403 n762__i1__i14__net1 n757__i1__i14__net1 22.45e-3
ri1405 n757__i1__i14__net1 n755__i1__i14__net1 18.86e-3
ri1407 n755__i1__i14__net1 n751__i1__i14__net1 22.45e-3
ri1409 n751__i1__i14__net1 n747__i1__i14__net1 18.86e-3
ri1411 n747__i1__i14__net1 n743__i1__i14__net1 21.86e-3
ri1413 n743__i1__i14__net1 n739__i1__i14__net1 18.86e-3
ri1415 n739__i1__i14__net1 n735__i1__i14__net1 22.45e-3
ri1417 n735__i1__i14__net1 n731__i1__i14__net1 18.86e-3
ri1419 n731__i1__i14__net1 n727__i1__i14__net1 22.45e-3
ri1421 n727__i1__i14__net1 n723__i1__i14__net1 18.86e-3
ri1423 n723__i1__i14__net1 n719__i1__i14__net1 22.45e-3
ri1425 n719__i1__i14__net1 n711__i1__i14__net1 18.86e-3
ri1427 n711__i1__i14__net1 n698__i1__i14__net1 22.45e-3
ri1429 n698__i1__i14__net1 n695__i1__i14__net1 18.86e-3
ri1431 n695__i1__i14__net1 n681__i1__i14__net1 22.45e-3
ri1433 n681__i1__i14__net1 n677__i1__i14__net1 18.86e-3
ri1435 n677__i1__i14__net1 n665__i1__i14__net1 22.45e-3
ri1437 n665__i1__i14__net1 n663__i1__i14__net1 18.86e-3
ri1439 n663__i1__i14__net1 n655__i1__i14__net1 22.45e-3
ri1441 n655__i1__i14__net1 n642__i1__i14__net1 18.86e-3
ri1443 n642__i1__i14__net1 n635__i1__i14__net1 21.86e-3
ri1445 n635__i1__i14__net1 n627__i1__i14__net1 18.86e-3
ri1447 n627__i1__i14__net1 n623__i1__i14__net1 22.45e-3
ri1449 n623__i1__i14__net1 n615__i1__i14__net1 18.86e-3
ri1451 n615__i1__i14__net1 n603__i1__i14__net1 22.45e-3
ri1453 n603__i1__i14__net1 n599__i1__i14__net1 18.86e-3
ri1455 n599__i1__i14__net1 n586__i1__i14__net1 22.45e-3
ri1457 n586__i1__i14__net1 n583__i1__i14__net1 18.86e-3
ri1459 n583__i1__i14__net1 n575__i1__i14__net1 22.45e-3
ri1461 n575__i1__i14__net1 n567__i1__i14__net1 18.86e-3
ri1463 n567__i1__i14__net1 n559__i1__i14__net1 22.45e-3
ri1465 n559__i1__i14__net1 n551__i1__i14__net1 18.86e-3
ri1467 n551__i1__i14__net1 n539__i1__i14__net1 21.86e-3
ri1469 n539__i1__i14__net1 n535__i1__i14__net1 18.86e-3
ri1471 n535__i1__i14__net1 n521__i1__i14__net1 22.45e-3
ri1473 n521__i1__i14__net1 n519__i1__i14__net1 18.86e-3
ri1475 n519__i1__i14__net1 n511__i1__i14__net1 22.45e-3
ri1477 n511__i1__i14__net1 n503__i1__i14__net1 18.86e-3
ri1479 n503__i1__i14__net1 n491__i1__i14__net1 22.45e-3
ri1481 n491__i1__i14__net1 n487__i1__i14__net1 18.86e-3
ri1483 n487__i1__i14__net1 n475__i1__i14__net1 22.45e-3
ri1485 n475__i1__i14__net1 n469__i1__i14__net1 18.86e-3
ri1487 n469__i1__i14__net1 n463__i1__i14__net1 22.45e-3
ri1489 n463__i1__i14__net1 n455__i1__i14__net1 18.86e-3
ri1491 n455__i1__i14__net1 n445__i1__i14__net1 22.45e-3
ri1493 n445__i1__i14__net1 n439__i1__i14__net1 18.86e-3
ri1495 n439__i1__i14__net1 n429__i1__i14__net1 22.45e-3
ri1497 n429__i1__i14__net1 n419__i1__i14__net1 18.86e-3
ri1499 n419__i1__i14__net1 n411__i1__i14__net1 23.05e-3
ri1501 n411__i1__i14__net1 n403__i1__i14__net1 18.86e-3
ri1503 n403__i1__i14__net1 n398__i1__i14__net1 22.45e-3
ri1505 n398__i1__i14__net1 n387__i1__i14__net1 18.86e-3
ri1507 n387__i1__i14__net1 n383__i1__i14__net1 23.05e-3
ri1509 n383__i1__i14__net1 n371__i1__i14__net1 18.86e-3
ri1511 n371__i1__i14__net1 n367__i1__i14__net1 22.45e-3
ri1513 n367__i1__i14__net1 n355__i1__i14__net1 18.86e-3
ri1515 n355__i1__i14__net1 n351__i1__i14__net1 22.45e-3
ri1517 n351__i1__i14__net1 n339__i1__i14__net1 18.86e-3
ri1519 n339__i1__i14__net1 n331__i1__i14__net1 22.45e-3
ri1521 n331__i1__i14__net1 n323__i1__i14__net1 18.86e-3
ri1523 n323__i1__i14__net1 n318__i1__i14__net1 21.86e-3
ri1525 n318__i1__i14__net1 n311__i1__i14__net1 18.86e-3
ri1527 n311__i1__i14__net1 n298__i1__i14__net1 22.45e-3
ri1529 n298__i1__i14__net1 n291__i1__i14__net1 18.86e-3
ri1531 n291__i1__i14__net1 n283__i1__i14__net1 22.45e-3
ri1533 n283__i1__i14__net1 n277__i1__i14__net1 18.86e-3
ri1535 n277__i1__i14__net1 n267__i1__i14__net1 22.45e-3
ri1537 n267__i1__i14__net1 n263__i1__i14__net1 18.86e-3
ri1539 n263__i1__i14__net1 n250__i1__i14__net1 22.45e-3
ri1541 n250__i1__i14__net1 n247__i1__i14__net1 18.86e-3
ri1543 n247__i1__i14__net1 n235__i1__i14__net1 22.45e-3
ri1545 n235__i1__i14__net1 n231__i1__i14__net1 18.86e-3
ri1547 n231__i1__i14__net1 n223__i1__i14__net1 22.45e-3
ri1549 n223__i1__i14__net1 n215__i1__i14__net1 18.86e-3
ri1551 n215__i1__i14__net1 n206__i1__i14__net1 22.45e-3
ri1553 n206__i1__i14__net1 n193__i1__i14__net1 18.86e-3
ri1555 n193__i1__i14__net1 n191__i1__i14__net1 21.86e-3
ri1557 n191__i1__i14__net1 n183__i1__i14__net1 18.86e-3
ri1559 n183__i1__i14__net1 n170__i1__i14__net1 22.45e-3
ri1561 n170__i1__i14__net1 n167__i1__i14__net1 18.86e-3
ri1563 n167__i1__i14__net1 n155__i1__i14__net1 22.45e-3
ri1565 n155__i1__i14__net1 n151__i1__i14__net1 18.86e-3
ri1567 n151__i1__i14__net1 n139__i1__i14__net1 22.45e-3
ri1569 n139__i1__i14__net1 n135__i1__i14__net1 18.86e-3
ri1571 n135__i1__i14__net1 n121__i1__i14__net1 22.45e-3
ri1573 n121__i1__i14__net1 n119__i1__i14__net1 18.86e-3
ri1575 n119__i1__i14__net1 n111__i1__i14__net1 22.45e-3
ri1577 n111__i1__i14__net1 n103__i1__i14__net1 18.86e-3
ri1579 n103__i1__i14__net1 n95__i1__i14__net1 21.86e-3
ri1581 n95__i1__i14__net1 n85__i1__i14__net1 18.86e-3
ri1583 n85__i1__i14__net1 n75__i1__i14__net1 22.45e-3
ri1585 n75__i1__i14__net1 n71__i1__i14__net1 18.86e-3
ri1587 n71__i1__i14__net1 n63__i1__i14__net1 25.1e-3
ri1589 n30__i5__i6__net31 n31__i5__i6__net31 500e-3
ri1590 n10__i5__i8__net1 n8__i5__i8__net1 250e-3
ri1591 n51__reset n52__reset 500e-3
ri1592 n36__shift n37__shift 500e-3
ri1593 n16__i5__i8__net2 n18__i5__i8__net2 250e-3
ri1594 n14__i5__r0 n15__i5__r0 166.7e-3
ri1595 n24__i5__i8__net1 n25__i5__i8__net1 500e-3
ri1596 n9__i5__i8__net5 n10__i5__i8__net5 250e-3
ri1597 n42__i5__i6__net31 n43__i5__i6__net31 500e-3
ri1598 n68__i5__clk_buf n66__i5__clk_buf 1.3551
ri1599 n66__i5__clk_buf n69__i5__clk_buf 2.3274
ri1600 n69__i5__clk_buf n52__i5__clk_buf 266.6e-3
ri1601 n52__i5__clk_buf n70__i5__clk_buf 452.5e-3
ri1602 n70__i5__clk_buf n43__i5__clk_buf 723.2e-3
ri1603 n69__i5__clk_buf n59__i5__clk_buf 1.0857
ri1604 n70__i5__clk_buf n71__i5__clk_buf 1.8735
ri1605 n71__i5__clk_buf n36__i5__clk_buf 1.0857
ri1606 n43__i5__clk_buf n57__i5__clk_buf 1.2155
ri1607 n57__i5__clk_buf n64__i5__clk_buf 1.3551
ri1608 n71__i5__clk_buf n27__i5__clk_buf 266.6e-3
ri1609 n27__i5__clk_buf n16__i5__clk_buf 2.1805
ri1610 n36__i5__i8__net2 n33__i5__i8__net2 1.8551
ri1611 n70__reset n72__reset 250e-3
ri1612 n71__reset n55__reset 2.4328
ri1614 n40__shift n41__shift 200e-3
ri1615 n12__i5__i8__net5 n19__i5__i8__net5 250e-3
ri1616 n98__i5__clk4 n99__i5__clk4 500e-3
ri1617 n18__piso_out n19__piso_out 125e-3
ri1618 n38__i5__i8__net2 n39__i5__i8__net2 500e-3
ri1619 piso_outinv n3__piso_outinv 250e-3
ri1620 n1300__i1__i14__net1 n1286__i1__i14__net1 82.23e-3
ri1621 n1286__i1__i14__net1 n1247__i1__i14__net1 82.23e-3
ri1622 n1247__i1__i14__net1 n1208__i1__i14__net1 82.23e-3
ri1623 n1208__i1__i14__net1 n1169__i1__i14__net1 82.23e-3
ri1624 n1169__i1__i14__net1 n1130__i1__i14__net1 82.23e-3
ri1625 n1130__i1__i14__net1 n1066__i1__i14__net1 82.23e-3
ri1626 n1066__i1__i14__net1 n1052__i1__i14__net1 82.23e-3
ri1627 n1052__i1__i14__net1 n1013__i1__i14__net1 79.87e-3
ri1628 n1013__i1__i14__net1 n974__i1__i14__net1 82.23e-3
ri1629 n974__i1__i14__net1 n935__i1__i14__net1 82.23e-3
ri1630 n935__i1__i14__net1 n896__i1__i14__net1 82.23e-3
ri1631 n896__i1__i14__net1 n857__i1__i14__net1 82.23e-3
ri1632 n857__i1__i14__net1 n818__i1__i14__net1 82.23e-3
ri1633 n818__i1__i14__net1 n779__i1__i14__net1 172.9e-3
ri1634 n1304__i1__i14__net1 n1288__i1__i14__net1 82.23e-3
ri1635 n1288__i1__i14__net1 n1249__i1__i14__net1 82.23e-3
ri1636 n1249__i1__i14__net1 n1210__i1__i14__net1 82.23e-3
ri1637 n1210__i1__i14__net1 n1171__i1__i14__net1 82.23e-3
ri1638 n1171__i1__i14__net1 n1132__i1__i14__net1 82.23e-3
ri1639 n1132__i1__i14__net1 n1070__i1__i14__net1 82.23e-3
ri1640 n1070__i1__i14__net1 n1054__i1__i14__net1 82.23e-3
ri1641 n1054__i1__i14__net1 n1015__i1__i14__net1 79.87e-3
ri1642 n1015__i1__i14__net1 n976__i1__i14__net1 82.23e-3
ri1643 n976__i1__i14__net1 n937__i1__i14__net1 82.23e-3
ri1644 n937__i1__i14__net1 n898__i1__i14__net1 82.23e-3
ri1645 n898__i1__i14__net1 n859__i1__i14__net1 82.23e-3
ri1646 n859__i1__i14__net1 n820__i1__i14__net1 82.23e-3
ri1647 n820__i1__i14__net1 n781__i1__i14__net1 172.9e-3
ri1648 n1299__i1__i14__net1 n1285__i1__i14__net1 82.59e-3
ri1649 n1285__i1__i14__net1 n1246__i1__i14__net1 82.59e-3
ri1650 n1246__i1__i14__net1 n1207__i1__i14__net1 82.59e-3
ri1651 n1207__i1__i14__net1 n1168__i1__i14__net1 82.59e-3
ri1652 n1168__i1__i14__net1 n1129__i1__i14__net1 82.59e-3
ri1653 n1129__i1__i14__net1 n1065__i1__i14__net1 82.59e-3
ri1654 n1065__i1__i14__net1 n1051__i1__i14__net1 82.59e-3
ri1655 n1051__i1__i14__net1 n1012__i1__i14__net1 80.23e-3
ri1656 n1012__i1__i14__net1 n973__i1__i14__net1 82.59e-3
ri1657 n973__i1__i14__net1 n934__i1__i14__net1 82.59e-3
ri1658 n934__i1__i14__net1 n895__i1__i14__net1 82.59e-3
ri1659 n895__i1__i14__net1 n856__i1__i14__net1 82.59e-3
ri1660 n856__i1__i14__net1 n817__i1__i14__net1 82.59e-3
ri1661 n817__i1__i14__net1 n778__i1__i14__net1 132e-3
ri1662 n1303__i1__i14__net1 n1287__i1__i14__net1 82.59e-3
ri1663 n1287__i1__i14__net1 n1248__i1__i14__net1 82.59e-3
ri1664 n1248__i1__i14__net1 n1209__i1__i14__net1 82.59e-3
ri1665 n1209__i1__i14__net1 n1170__i1__i14__net1 82.59e-3
ri1666 n1170__i1__i14__net1 n1131__i1__i14__net1 82.59e-3
ri1667 n1131__i1__i14__net1 n1069__i1__i14__net1 82.59e-3
ri1668 n1069__i1__i14__net1 n1053__i1__i14__net1 82.59e-3
ri1669 n1053__i1__i14__net1 n1014__i1__i14__net1 80.23e-3
ri1670 n1014__i1__i14__net1 n975__i1__i14__net1 82.59e-3
ri1671 n975__i1__i14__net1 n936__i1__i14__net1 82.59e-3
ri1672 n936__i1__i14__net1 n897__i1__i14__net1 82.59e-3
ri1673 n897__i1__i14__net1 n858__i1__i14__net1 82.59e-3
ri1674 n858__i1__i14__net1 n819__i1__i14__net1 82.59e-3
ri1675 n819__i1__i14__net1 n780__i1__i14__net1 173.1e-3
ri1676 n1307__i1__i14__net1 n1289__i1__i14__net1 82.59e-3
ri1677 n1289__i1__i14__net1 n1250__i1__i14__net1 82.59e-3
ri1678 n1250__i1__i14__net1 n1211__i1__i14__net1 82.59e-3
ri1679 n1211__i1__i14__net1 n1172__i1__i14__net1 82.59e-3
ri1680 n1172__i1__i14__net1 n1133__i1__i14__net1 82.59e-3
ri1681 n1133__i1__i14__net1 n1073__i1__i14__net1 82.59e-3
ri1682 n1073__i1__i14__net1 n1055__i1__i14__net1 82.59e-3
ri1683 n1055__i1__i14__net1 n1016__i1__i14__net1 80.23e-3
ri1684 n1016__i1__i14__net1 n977__i1__i14__net1 82.59e-3
ri1685 n977__i1__i14__net1 n938__i1__i14__net1 82.59e-3
ri1686 n938__i1__i14__net1 n899__i1__i14__net1 82.59e-3
ri1687 n899__i1__i14__net1 n860__i1__i14__net1 82.59e-3
ri1688 n860__i1__i14__net1 n821__i1__i14__net1 82.59e-3
ri1689 n821__i1__i14__net1 n782__i1__i14__net1 173.1e-3
ri1690 n1308__i1__i14__net1 n1290__i1__i14__net1 82.59e-3
ri1691 n1290__i1__i14__net1 n1251__i1__i14__net1 82.59e-3
ri1692 n1251__i1__i14__net1 n1212__i1__i14__net1 82.59e-3
ri1693 n1212__i1__i14__net1 n1173__i1__i14__net1 82.59e-3
ri1694 n1173__i1__i14__net1 n1134__i1__i14__net1 82.59e-3
ri1695 n1134__i1__i14__net1 n1074__i1__i14__net1 82.59e-3
ri1696 n1074__i1__i14__net1 n1056__i1__i14__net1 82.59e-3
ri1697 n1056__i1__i14__net1 n1017__i1__i14__net1 80.23e-3
ri1698 n1017__i1__i14__net1 n978__i1__i14__net1 82.59e-3
ri1699 n978__i1__i14__net1 n939__i1__i14__net1 82.59e-3
ri1700 n939__i1__i14__net1 n900__i1__i14__net1 82.59e-3
ri1701 n900__i1__i14__net1 n861__i1__i14__net1 82.59e-3
ri1702 n861__i1__i14__net1 n822__i1__i14__net1 82.59e-3
ri1703 n822__i1__i14__net1 n783__i1__i14__net1 173.7e-3
ri1704 n1311__i1__i14__net1 n1291__i1__i14__net1 82.59e-3
ri1705 n1291__i1__i14__net1 n1252__i1__i14__net1 82.59e-3
ri1706 n1252__i1__i14__net1 n1213__i1__i14__net1 82.59e-3
ri1707 n1213__i1__i14__net1 n1174__i1__i14__net1 82.59e-3
ri1708 n1174__i1__i14__net1 n1135__i1__i14__net1 82.59e-3
ri1709 n1135__i1__i14__net1 n1077__i1__i14__net1 82.59e-3
ri1710 n1077__i1__i14__net1 n1057__i1__i14__net1 82.59e-3
ri1711 n1057__i1__i14__net1 n1018__i1__i14__net1 80.23e-3
ri1712 n1018__i1__i14__net1 n979__i1__i14__net1 82.59e-3
ri1713 n979__i1__i14__net1 n940__i1__i14__net1 82.59e-3
ri1714 n940__i1__i14__net1 n901__i1__i14__net1 82.59e-3
ri1715 n901__i1__i14__net1 n862__i1__i14__net1 82.59e-3
ri1716 n862__i1__i14__net1 n823__i1__i14__net1 82.59e-3
ri1717 n823__i1__i14__net1 n784__i1__i14__net1 173.1e-3
ri1718 n1312__i1__i14__net1 n1292__i1__i14__net1 82.59e-3
ri1719 n1292__i1__i14__net1 n1253__i1__i14__net1 82.59e-3
ri1720 n1253__i1__i14__net1 n1214__i1__i14__net1 82.59e-3
ri1721 n1214__i1__i14__net1 n1175__i1__i14__net1 82.59e-3
ri1722 n1175__i1__i14__net1 n1136__i1__i14__net1 82.59e-3
ri1723 n1136__i1__i14__net1 n1078__i1__i14__net1 82.59e-3
ri1724 n1078__i1__i14__net1 n1058__i1__i14__net1 82.59e-3
ri1725 n1058__i1__i14__net1 n1019__i1__i14__net1 80.23e-3
ri1726 n1019__i1__i14__net1 n980__i1__i14__net1 82.59e-3
ri1727 n980__i1__i14__net1 n941__i1__i14__net1 82.59e-3
ri1728 n941__i1__i14__net1 n902__i1__i14__net1 82.59e-3
ri1729 n902__i1__i14__net1 n863__i1__i14__net1 82.59e-3
ri1730 n863__i1__i14__net1 n824__i1__i14__net1 82.59e-3
ri1731 n824__i1__i14__net1 n785__i1__i14__net1 173.7e-3
ri1732 n1315__i1__i14__net1 n1293__i1__i14__net1 82.59e-3
ri1733 n1293__i1__i14__net1 n1254__i1__i14__net1 82.59e-3
ri1734 n1254__i1__i14__net1 n1215__i1__i14__net1 82.59e-3
ri1735 n1215__i1__i14__net1 n1176__i1__i14__net1 82.59e-3
ri1736 n1176__i1__i14__net1 n1137__i1__i14__net1 82.59e-3
ri1737 n1137__i1__i14__net1 n1081__i1__i14__net1 82.59e-3
ri1738 n1081__i1__i14__net1 n1059__i1__i14__net1 82.59e-3
ri1739 n1059__i1__i14__net1 n1020__i1__i14__net1 80.23e-3
ri1740 n1020__i1__i14__net1 n981__i1__i14__net1 82.59e-3
ri1741 n981__i1__i14__net1 n942__i1__i14__net1 82.59e-3
ri1742 n942__i1__i14__net1 n903__i1__i14__net1 82.59e-3
ri1743 n903__i1__i14__net1 n864__i1__i14__net1 82.59e-3
ri1744 n864__i1__i14__net1 n825__i1__i14__net1 82.59e-3
ri1745 n825__i1__i14__net1 n786__i1__i14__net1 173.1e-3
ri1746 n1316__i1__i14__net1 n1294__i1__i14__net1 82.59e-3
ri1747 n1294__i1__i14__net1 n1255__i1__i14__net1 82.59e-3
ri1748 n1255__i1__i14__net1 n1216__i1__i14__net1 82.59e-3
ri1749 n1216__i1__i14__net1 n1177__i1__i14__net1 82.59e-3
ri1750 n1177__i1__i14__net1 n1138__i1__i14__net1 82.59e-3
ri1751 n1138__i1__i14__net1 n1082__i1__i14__net1 82.59e-3
ri1752 n1082__i1__i14__net1 n1060__i1__i14__net1 82.59e-3
ri1753 n1060__i1__i14__net1 n1021__i1__i14__net1 80.23e-3
ri1754 n1021__i1__i14__net1 n982__i1__i14__net1 82.59e-3
ri1755 n982__i1__i14__net1 n943__i1__i14__net1 82.59e-3
ri1756 n943__i1__i14__net1 n904__i1__i14__net1 82.59e-3
ri1757 n904__i1__i14__net1 n865__i1__i14__net1 82.59e-3
ri1758 n865__i1__i14__net1 n826__i1__i14__net1 82.59e-3
ri1759 n826__i1__i14__net1 n787__i1__i14__net1 173.1e-3
ri1760 n1319__i1__i14__net1 n1295__i1__i14__net1 82.59e-3
ri1761 n1295__i1__i14__net1 n1256__i1__i14__net1 82.59e-3
ri1762 n1256__i1__i14__net1 n1217__i1__i14__net1 82.59e-3
ri1763 n1217__i1__i14__net1 n1178__i1__i14__net1 82.59e-3
ri1764 n1178__i1__i14__net1 n1139__i1__i14__net1 82.59e-3
ri1765 n1139__i1__i14__net1 n1085__i1__i14__net1 82.59e-3
ri1766 n1085__i1__i14__net1 n1061__i1__i14__net1 82.59e-3
ri1767 n1061__i1__i14__net1 n1022__i1__i14__net1 80.23e-3
ri1768 n1022__i1__i14__net1 n983__i1__i14__net1 82.59e-3
ri1769 n983__i1__i14__net1 n944__i1__i14__net1 82.59e-3
ri1770 n944__i1__i14__net1 n905__i1__i14__net1 82.59e-3
ri1771 n905__i1__i14__net1 n866__i1__i14__net1 82.59e-3
ri1772 n866__i1__i14__net1 n827__i1__i14__net1 82.59e-3
ri1773 n827__i1__i14__net1 n788__i1__i14__net1 173.1e-3
ri1774 n1320__i1__i14__net1 n1296__i1__i14__net1 82.59e-3
ri1775 n1296__i1__i14__net1 n1257__i1__i14__net1 82.59e-3
ri1776 n1257__i1__i14__net1 n1218__i1__i14__net1 82.59e-3
ri1777 n1218__i1__i14__net1 n1179__i1__i14__net1 82.59e-3
ri1778 n1179__i1__i14__net1 n1140__i1__i14__net1 82.59e-3
ri1779 n1140__i1__i14__net1 n1086__i1__i14__net1 82.59e-3
ri1780 n1086__i1__i14__net1 n1062__i1__i14__net1 82.59e-3
ri1781 n1062__i1__i14__net1 n1023__i1__i14__net1 80.23e-3
ri1782 n1023__i1__i14__net1 n984__i1__i14__net1 82.59e-3
ri1783 n984__i1__i14__net1 n945__i1__i14__net1 82.59e-3
ri1784 n945__i1__i14__net1 n906__i1__i14__net1 82.59e-3
ri1785 n906__i1__i14__net1 n867__i1__i14__net1 82.59e-3
ri1786 n867__i1__i14__net1 n828__i1__i14__net1 82.59e-3
ri1787 n828__i1__i14__net1 n789__i1__i14__net1 173.1e-3
ri1788 n1323__i1__i14__net1 n1297__i1__i14__net1 82.59e-3
ri1789 n1297__i1__i14__net1 n1258__i1__i14__net1 82.59e-3
ri1790 n1258__i1__i14__net1 n1219__i1__i14__net1 82.59e-3
ri1791 n1219__i1__i14__net1 n1180__i1__i14__net1 82.59e-3
ri1792 n1180__i1__i14__net1 n1141__i1__i14__net1 82.59e-3
ri1793 n1141__i1__i14__net1 n1089__i1__i14__net1 82.59e-3
ri1794 n1089__i1__i14__net1 n1063__i1__i14__net1 82.59e-3
ri1795 n1063__i1__i14__net1 n1024__i1__i14__net1 80.23e-3
ri1796 n1024__i1__i14__net1 n985__i1__i14__net1 82.59e-3
ri1797 n985__i1__i14__net1 n946__i1__i14__net1 82.59e-3
ri1798 n946__i1__i14__net1 n907__i1__i14__net1 82.59e-3
ri1799 n907__i1__i14__net1 n868__i1__i14__net1 82.59e-3
ri1800 n868__i1__i14__net1 n829__i1__i14__net1 82.59e-3
ri1801 n829__i1__i14__net1 n790__i1__i14__net1 131.5e-3
ri1802 n1493__vddio n1472__vddio 82.59e-3
ri1803 n1472__vddio n1465__vddio 82.59e-3
ri1804 n1465__vddio n1444__vddio 82.59e-3
ri1805 n1444__vddio n1423__vddio 82.59e-3
ri1806 n1423__vddio n1392__vddio 82.59e-3
ri1807 n1392__vddio n1371__vddio 82.59e-3
ri1808 n1371__vddio n1337__vddio 82.59e-3
ri1809 n1337__vddio n1329__vddio 80.23e-3
ri1810 n1329__vddio n1308__vddio 82.59e-3
ri1811 n1308__vddio n1277__vddio 82.59e-3
ri1812 n1277__vddio n1242__vddio 82.59e-3
ri1813 n1242__vddio n1235__vddio 82.59e-3
ri1814 n1235__vddio n1214__vddio 82.59e-3
ri1815 n1214__vddio n1187__vddio 82.59e-3
ri1816 n1496__vddio n1475__vddio 82.59e-3
ri1817 n1475__vddio n1466__vddio 82.59e-3
ri1818 n1466__vddio n1445__vddio 82.59e-3
ri1819 n1445__vddio n1424__vddio 82.59e-3
ri1820 n1424__vddio n1393__vddio 82.59e-3
ri1821 n1393__vddio n1372__vddio 82.59e-3
ri1822 n1372__vddio n1338__vddio 82.59e-3
ri1823 n1338__vddio n1330__vddio 80.23e-3
ri1824 n1330__vddio n1309__vddio 82.59e-3
ri1825 n1309__vddio n1278__vddio 82.59e-3
ri1826 n1278__vddio n1245__vddio 82.59e-3
ri1827 n1245__vddio n1236__vddio 82.59e-3
ri1828 n1236__vddio n1215__vddio 82.59e-3
ri1829 n1215__vddio n1188__vddio 82.59e-3
ri1830 n1497__vddio n1476__vddio 82.59e-3
ri1831 n1476__vddio n1467__vddio 82.59e-3
ri1832 n1467__vddio n1446__vddio 82.59e-3
ri1833 n1446__vddio n1425__vddio 82.59e-3
ri1834 n1425__vddio n1394__vddio 82.59e-3
ri1835 n1394__vddio n1373__vddio 82.59e-3
ri1836 n1373__vddio n1341__vddio 82.59e-3
ri1837 n1341__vddio n1331__vddio 80.23e-3
ri1838 n1331__vddio n1310__vddio 82.59e-3
ri1839 n1310__vddio n1279__vddio 82.59e-3
ri1840 n1279__vddio n1246__vddio 82.59e-3
ri1841 n1246__vddio n1237__vddio 82.59e-3
ri1842 n1237__vddio n1216__vddio 82.59e-3
ri1843 n1216__vddio n1189__vddio 82.59e-3
ri1844 n1500__vddio n1479__vddio 82.59e-3
ri1845 n1479__vddio n1468__vddio 82.59e-3
ri1846 n1468__vddio n1447__vddio 82.59e-3
ri1847 n1447__vddio n1426__vddio 82.59e-3
ri1848 n1426__vddio n1395__vddio 82.59e-3
ri1849 n1395__vddio n1374__vddio 82.59e-3
ri1850 n1374__vddio n1342__vddio 82.59e-3
ri1851 n1342__vddio n1332__vddio 80.23e-3
ri1852 n1332__vddio n1311__vddio 82.59e-3
ri1853 n1311__vddio n1280__vddio 82.59e-3
ri1854 n1280__vddio n1249__vddio 82.59e-3
ri1855 n1249__vddio n1238__vddio 82.59e-3
ri1856 n1238__vddio n1217__vddio 82.59e-3
ri1857 n1217__vddio n1190__vddio 82.59e-3
ri1858 n1501__vddio n1480__vddio 82.59e-3
ri1859 n1480__vddio n1469__vddio 82.59e-3
ri1860 n1469__vddio n1448__vddio 82.59e-3
ri1861 n1448__vddio n1427__vddio 82.59e-3
ri1862 n1427__vddio n1396__vddio 82.59e-3
ri1863 n1396__vddio n1375__vddio 82.59e-3
ri1864 n1375__vddio n1345__vddio 82.59e-3
ri1865 n1345__vddio n1333__vddio 80.23e-3
ri1866 n1333__vddio n1312__vddio 82.59e-3
ri1867 n1312__vddio n1281__vddio 82.59e-3
ri1868 n1281__vddio n1250__vddio 82.59e-3
ri1869 n1250__vddio n1239__vddio 82.59e-3
ri1870 n1239__vddio n1218__vddio 82.59e-3
ri1871 n1218__vddio n1191__vddio 82.59e-3
ri1872 n1504__vddio n1483__vddio 82.59e-3
ri1873 n1483__vddio n1470__vddio 82.59e-3
ri1874 n1470__vddio n1449__vddio 82.59e-3
ri1875 n1449__vddio n1428__vddio 82.59e-3
ri1876 n1428__vddio n1397__vddio 82.59e-3
ri1877 n1397__vddio n1376__vddio 82.59e-3
ri1878 n1376__vddio n1346__vddio 82.59e-3
ri1879 n1346__vddio n1334__vddio 80.23e-3
ri1880 n1334__vddio n1313__vddio 82.59e-3
ri1881 n1313__vddio n1282__vddio 82.59e-3
ri1882 n1282__vddio n1253__vddio 82.59e-3
ri1883 n1253__vddio n1240__vddio 82.59e-3
ri1884 n1240__vddio n1219__vddio 82.59e-3
ri1885 n1219__vddio n1192__vddio 82.59e-3
ri1886 n1505__vddio n1484__vddio 82.59e-3
ri1887 n1484__vddio n1471__vddio 82.59e-3
ri1888 n1471__vddio n1450__vddio 82.59e-3
ri1889 n1450__vddio n1429__vddio 82.59e-3
ri1890 n1429__vddio n1398__vddio 82.59e-3
ri1891 n1398__vddio n1377__vddio 82.59e-3
ri1892 n1377__vddio n1349__vddio 82.59e-3
ri1893 n1349__vddio n1335__vddio 80.23e-3
ri1894 n1335__vddio n1314__vddio 82.59e-3
ri1895 n1314__vddio n1283__vddio 82.59e-3
ri1896 n1283__vddio n1254__vddio 82.59e-3
ri1897 n1254__vddio n1241__vddio 82.59e-3
ri1898 n1241__vddio n1220__vddio 82.59e-3
ri1899 n1220__vddio n1193__vddio 82.59e-3
ri1900 n1507__vddio n1508__vddio 165.9e-3
ri1901 n1508__vddio n1509__vddio 82.59e-3
ri1902 n1509__vddio n1510__vddio 82.59e-3
ri1903 n1510__vddio n1511__vddio 82.59e-3
ri1904 n1511__vddio n1512__vddio 82.59e-3
ri1905 n1512__vddio n1513__vddio 82.59e-3
ri1906 n1513__vddio n1514__vddio 82.59e-3
ri1907 n1514__vddio n1515__vddio 80.23e-3
ri1908 n1515__vddio n1516__vddio 82.59e-3
ri1909 n1516__vddio n1517__vddio 82.59e-3
ri1910 n1517__vddio n1518__vddio 82.59e-3
ri1911 n1518__vddio n1519__vddio 82.59e-3
ri1912 n1519__vddio n1520__vddio 82.59e-3
ri1913 n1520__vddio n1186__vddio 165.9e-3
ri1914 n893__vss n894__vss 165.9e-3
ri1915 n894__vss n895__vss 82.59e-3
ri1916 n895__vss n896__vss 82.59e-3
ri1917 n896__vss n897__vss 82.59e-3
ri1918 n897__vss n898__vss 82.59e-3
ri1919 n898__vss n899__vss 82.59e-3
ri1920 n899__vss n900__vss 82.59e-3
ri1921 n900__vss n901__vss 80.23e-3
ri1922 n901__vss n902__vss 82.59e-3
ri1923 n902__vss n903__vss 82.59e-3
ri1924 n903__vss n904__vss 82.59e-3
ri1925 n904__vss n905__vss 82.59e-3
ri1926 n905__vss n906__vss 82.59e-3
ri1927 n906__vss n711__vss 165.9e-3
ri1928 n885__vss n872__vss 82.59e-3
ri1929 n872__vss n868__vss 82.59e-3
ri1930 n868__vss n855__vss 82.59e-3
ri1931 n855__vss n842__vss 82.59e-3
ri1932 n842__vss n829__vss 82.59e-3
ri1933 n829__vss n816__vss 82.59e-3
ri1934 n816__vss n795__vss 82.59e-3
ri1935 n795__vss n790__vss 80.23e-3
ri1936 n790__vss n777__vss 82.59e-3
ri1937 n777__vss n764__vss 82.59e-3
ri1938 n764__vss n742__vss 82.59e-3
ri1939 n742__vss n738__vss 82.59e-3
ri1940 n738__vss n725__vss 82.59e-3
ri1941 n725__vss n712__vss 82.59e-3
ri1942 n888__vss n875__vss 82.59e-3
ri1943 n875__vss n869__vss 82.59e-3
ri1944 n869__vss n856__vss 82.59e-3
ri1945 n856__vss n843__vss 82.59e-3
ri1946 n843__vss n830__vss 82.59e-3
ri1947 n830__vss n817__vss 82.59e-3
ri1948 n817__vss n796__vss 82.59e-3
ri1949 n796__vss n791__vss 80.23e-3
ri1950 n791__vss n778__vss 82.59e-3
ri1951 n778__vss n765__vss 82.59e-3
ri1952 n765__vss n745__vss 82.59e-3
ri1953 n745__vss n739__vss 82.59e-3
ri1954 n739__vss n726__vss 82.59e-3
ri1955 n726__vss n713__vss 82.59e-3
ri1956 n889__vss n876__vss 82.59e-3
ri1957 n876__vss n870__vss 82.59e-3
ri1958 n870__vss n857__vss 82.59e-3
ri1959 n857__vss n844__vss 82.59e-3
ri1960 n844__vss n831__vss 82.59e-3
ri1961 n831__vss n818__vss 82.59e-3
ri1962 n818__vss n799__vss 82.59e-3
ri1963 n799__vss n792__vss 80.23e-3
ri1964 n792__vss n779__vss 82.59e-3
ri1965 n779__vss n766__vss 82.59e-3
ri1966 n766__vss n746__vss 82.59e-3
ri1967 n746__vss n740__vss 82.59e-3
ri1968 n740__vss n727__vss 82.59e-3
ri1969 n727__vss n714__vss 82.59e-3
ri1970 n892__vss n879__vss 82.59e-3
ri1971 n879__vss n871__vss 82.59e-3
ri1972 n871__vss n858__vss 82.59e-3
ri1973 n858__vss n845__vss 82.59e-3
ri1974 n845__vss n832__vss 82.59e-3
ri1975 n832__vss n819__vss 82.59e-3
ri1976 n819__vss n800__vss 82.59e-3
ri1977 n800__vss n793__vss 80.23e-3
ri1978 n793__vss n780__vss 82.59e-3
ri1979 n780__vss n767__vss 82.59e-3
ri1980 n767__vss n749__vss 82.59e-3
ri1981 n749__vss n741__vss 82.59e-3
ri1982 n741__vss n728__vss 82.59e-3
ri1983 n728__vss n715__vss 82.59e-3
ri1985 n385__vdd n387__vdd 447.8e-3
ri1987 n387__vdd n389__vdd 447.8e-3
ri1989 n389__vdd n391__vdd 447.8e-3
ri1991 n391__vdd n393__vdd 447.8e-3
ri1992 n393__vdd n384__vdd 12.5e-3
ri1993 n376__vdd n385__vdd 12.5e-3
ri1994 n378__vdd n387__vdd 12.5e-3
ri1995 n380__vdd n389__vdd 12.5e-3
ri1996 n382__vdd n391__vdd 12.5e-3
ri1998 n223__i1__net2 n225__i1__net2 384.5e-3
ri1999 n225__i1__net2 n226__i1__net2 91.38e-3
ri2000 n226__i1__net2 n227__i1__net2 90.6e-3
ri2001 n227__i1__net2 n228__i1__net2 182e-3
ri2002 n228__i1__net2 n229__i1__net2 154.7e-3
ri2003 n223__i1__net2 n219__i1__net2 18.97e-3
ri2005 n219__i1__net2 n213__i1__net2 22.52e-3
ri2007 n213__i1__net2 n211__i1__net2 18.97e-3
ri2009 n211__i1__net2 n207__i1__net2 22.52e-3
ri2011 n207__i1__net2 n203__i1__net2 18.97e-3
ri2013 n203__i1__net2 n199__i1__net2 22.52e-3
ri2015 n199__i1__net2 n195__i1__net2 18.97e-3
ri2017 n195__i1__net2 n191__i1__net2 21.93e-3
ri2019 n191__i1__net2 n186__i1__net2 18.97e-3
ri2021 n186__i1__net2 n179__i1__net2 22.52e-3
ri2023 n179__i1__net2 n175__i1__net2 18.97e-3
ri2025 n175__i1__net2 n173__i1__net2 22.52e-3
ri2027 n173__i1__net2 n165__i1__net2 18.97e-3
ri2029 n165__i1__net2 n161__i1__net2 22.52e-3
ri2031 n161__i1__net2 n159__i1__net2 18.97e-3
ri2033 n159__i1__net2 n151__i1__net2 22.52e-3
ri2035 n151__i1__net2 n143__i1__net2 18.97e-3
ri2037 n143__i1__net2 n131__i1__net2 22.52e-3
ri2039 n131__i1__net2 n125__i1__net2 18.97e-3
ri2041 n125__i1__net2 n117__i1__net2 22.52e-3
ri2043 n117__i1__net2 n111__i1__net2 18.97e-3
ri2045 n111__i1__net2 n99__i1__net2 22.52e-3
ri2047 n99__i1__net2 n91__i1__net2 18.97e-3
ri2049 n91__i1__net2 n82__i1__net2 21.93e-3
ri2051 n82__i1__net2 n79__i1__net2 18.97e-3
ri2053 n79__i1__net2 n71__i1__net2 22.52e-3
ri2055 n71__i1__net2 n63__i1__net2 18.97e-3
ri2057 n57__i1__i12__net1 n58__i1__i12__net1 175.8e-3
ri2058 n58__i1__i12__net1 n59__i1__i12__net1 105.9e-3
ri2059 n59__i1__i12__net1 n39__i1__i12__net1 91.22e-3
ri2060 n39__i1__i12__net1 n40__i1__i12__net1 108.8e-3
ri2061 n40__i1__i12__net1 n36__i1__i12__net1 47.91e-3
ri2062 n36__i1__i12__net1 n35__i1__i12__net1 178.2e-3
ri2063 n35__i1__i12__net1 n60__i1__i12__net1 62.94e-3
ri2064 n60__i1__i12__net1 n32__i1__i12__net1 75.16e-3
ri2065 n58__i1__i12__net1 n52__i1__i12__net1 32.85e-3
ri2067 n58__i1__i12__net1 n51__i1__i12__net1 40.41e-3
ri2069 n59__i1__i12__net1 n44__i1__i12__net1 32.78e-3
ri2071 n59__i1__i12__net1 n43__i1__i12__net1 39.87e-3
ri2073 n35__i1__i12__net1 n39__i1__i12__net1 26.15e-3
ri2074 n60__i1__i12__net1 n31__i1__i12__net1 81.63e-3
ri2075 n21__i1__net4 n19__i1__net4 146.5e-3
ri2077 n19__i1__net4 n15__i1__net4 17.28e-3
ri2080 n1734__vddio n1736__vddio 212.2e-3
ri2081 n1736__vddio n1737__vddio 8.333e-3
ri2082 n1730__vddio n1734__vddio 16.67e-3
ri2083 n1732__vddio n1736__vddio 8.333e-3
ri2084 n29__piso_out n30__piso_out 250e-3
ri2085 n18__piso_outinv n19__piso_outinv 250e-3
ri2086 n202__i1__i13__net1 n205__i1__i13__net1 117.8e-3
ri2087 n205__i1__i13__net1 n215__i1__i13__net1 82.3e-3
ri2088 n215__i1__i13__net1 n216__i1__i13__net1 85.36e-3
ri2089 n216__i1__i13__net1 n217__i1__i13__net1 90.43e-3
ri2090 n217__i1__i13__net1 n218__i1__i13__net1 102.2e-3
ri2091 n218__i1__i13__net1 n219__i1__i13__net1 102.2e-3
ri2092 n219__i1__i13__net1 n220__i1__i13__net1 102.2e-3
ri2093 n220__i1__i13__net1 n221__i1__i13__net1 102.2e-3
ri2094 n221__i1__i13__net1 n222__i1__i13__net1 102.2e-3
ri2095 n222__i1__i13__net1 n223__i1__i13__net1 102.2e-3
ri2096 n223__i1__i13__net1 n224__i1__i13__net1 103e-3
ri2097 n224__i1__i13__net1 n225__i1__i13__net1 103e-3
ri2098 n225__i1__i13__net1 n226__i1__i13__net1 77.03e-3
ri2099 n226__i1__i13__net1 n64__i1__i13__net1 29.56e-3
ri2101 n215__i1__i13__net1 n206__i1__i13__net1 147.7e-3
ri2102 n206__i1__i13__net1 n209__i1__i13__net1 113.6e-3
ri2103 n209__i1__i13__net1 n212__i1__i13__net1 119.2e-3
ri2104 n216__i1__i13__net1 n201__i1__i13__net1 41.61e-3
ri2105 n216__i1__i13__net1 n200__i1__i13__net1 42.95e-3
ri2106 n217__i1__i13__net1 n197__i1__i13__net1 28.84e-3
ri2108 n217__i1__i13__net1 n196__i1__i13__net1 29.76e-3
ri2110 n218__i1__i13__net1 n193__i1__i13__net1 28.84e-3
ri2112 n218__i1__i13__net1 n192__i1__i13__net1 29.76e-3
ri2114 n219__i1__i13__net1 n144__i1__i13__net1 28.84e-3
ri2116 n219__i1__i13__net1 n143__i1__i13__net1 29.76e-3
ri2118 n220__i1__i13__net1 n136__i1__i13__net1 28.84e-3
ri2120 n220__i1__i13__net1 n135__i1__i13__net1 29.76e-3
ri2122 n221__i1__i13__net1 n128__i1__i13__net1 28.84e-3
ri2124 n221__i1__i13__net1 n127__i1__i13__net1 29.76e-3
ri2126 n222__i1__i13__net1 n116__i1__i13__net1 28.84e-3
ri2128 n222__i1__i13__net1 n115__i1__i13__net1 29.76e-3
ri2130 n223__i1__i13__net1 n108__i1__i13__net1 28.84e-3
ri2132 n223__i1__i13__net1 n105__i1__i13__net1 29.76e-3
ri2134 n224__i1__i13__net1 n96__i1__i13__net1 28.34e-3
ri2136 n224__i1__i13__net1 n93__i1__i13__net1 29.25e-3
ri2138 n225__i1__i13__net1 n76__i1__i13__net1 28.84e-3
ri2140 n225__i1__i13__net1 n75__i1__i13__net1 29.76e-3
ri2142 n226__i1__i13__net1 n63__i1__i13__net1 30.48e-3
ri2144 n1714__vss n1715__vss 69.76e-3
ri2145 n1715__vss n1716__vss 199.7e-3
ri2146 n1716__vss n1717__vss 2.406e-3
ri2147 n1717__vss n1718__vss 267e-3
ri2148 n1718__vss n1719__vss 2.406e-3
ri2149 n1719__vss n1720__vss 267e-3
ri2150 n1720__vss n1721__vss 2.406e-3
ri2151 n1721__vss n1722__vss 267e-3
ri2152 n1722__vss n1723__vss 2.406e-3
ri2153 n1723__vss n1724__vss 267e-3
ri2154 n1724__vss n1725__vss 2.406e-3
ri2155 n1725__vss n1726__vss 267e-3
ri2156 n1726__vss n1727__vss 2.406e-3
ri2157 n1727__vss n1728__vss 267e-3
ri2158 n1728__vss n1729__vss 2.406e-3
ri2159 n1729__vss n1730__vss 267e-3
ri2160 n1730__vss n1731__vss 2.406e-3
ri2161 n1731__vss n1732__vss 267e-3
ri2162 n1732__vss n1733__vss 2.406e-3
ri2163 n1733__vss n1734__vss 267e-3
ri2164 n1734__vss n1735__vss 2.406e-3
ri2165 n1735__vss n1736__vss 267e-3
ri2166 n1736__vss n1737__vss 2.406e-3
ri2167 n1737__vss n1738__vss 267e-3
ri2168 n1738__vss n1739__vss 2.406e-3
ri2169 n1739__vss n1740__vss 267e-3
ri2170 n1740__vss n1741__vss 2.406e-3
ri2171 n1741__vss n1742__vss 267e-3
ri2172 n1742__vss n1743__vss 2.406e-3
ri2173 n1743__vss n1744__vss 267e-3
ri2174 n1744__vss n1745__vss 2.406e-3
ri2175 n1745__vss n1746__vss 267e-3
ri2176 n1746__vss n1010__vss 10.74e-3
ri2177 n1714__vss n1747__vss 212.2e-3
ri2178 n1747__vss n1748__vss 44.46e-3
ri2179 n1748__vss n1749__vss 224.7e-3
ri2180 n1749__vss n1750__vss 264.4e-3
ri2181 n1750__vss n1751__vss 157.3e-3
ri2182 n1751__vss n1752__vss 419.8e-3
ri2183 n1752__vss n1753__vss 277.2e-3
ri2184 n1753__vss n1713__vss 298.3e-3
ri2191 n1713__vss n1687__vss 3.012e-3
ri2205 n1687__vss n1675__vss 125e-3
ri2206 n1425__vss n1714__vss 8.333e-3
ri2207 n913__vss n1715__vss 16.67e-3
ri2208 n1427__vss n1716__vss 8.333e-3
ri2209 n919__vss n1717__vss 8.333e-3
ri2210 n1429__vss n1718__vss 8.333e-3
ri2211 n926__vss n1719__vss 8.333e-3
ri2212 n1431__vss n1720__vss 8.333e-3
ri2213 n934__vss n1721__vss 8.333e-3
ri2214 n1433__vss n1722__vss 8.333e-3
ri2215 n939__vss n1723__vss 8.333e-3
ri2216 n1435__vss n1724__vss 8.333e-3
ri2217 n944__vss n1725__vss 8.333e-3
ri2218 n1437__vss n1726__vss 8.333e-3
ri2219 n949__vss n1727__vss 8.333e-3
ri2220 n1439__vss n1728__vss 8.333e-3
ri2221 n954__vss n1729__vss 8.333e-3
ri2222 n1441__vss n1730__vss 8.333e-3
ri2223 n960__vss n1731__vss 8.333e-3
ri2224 n1443__vss n1732__vss 8.333e-3
ri2225 n966__vss n1733__vss 8.333e-3
ri2226 n1445__vss n1734__vss 8.333e-3
ri2227 n971__vss n1735__vss 8.333e-3
ri2228 n1447__vss n1736__vss 8.333e-3
ri2229 n978__vss n1737__vss 8.333e-3
ri2230 n1449__vss n1738__vss 8.333e-3
ri2231 n986__vss n1739__vss 8.333e-3
ri2232 n1451__vss n1740__vss 8.333e-3
ri2233 n991__vss n1741__vss 8.333e-3
ri2234 n1453__vss n1742__vss 8.333e-3
ri2235 n997__vss n1743__vss 8.333e-3
ri2236 n1455__vss n1744__vss 8.333e-3
ri2237 n1004__vss n1745__vss 8.333e-3
ri2238 n1457__vss n1746__vss 8.333e-3
ri2239 n1423__vss n1747__vss 16.67e-3
ri2240 n1586__vss n1748__vss 12.5e-3
ri2241 n1584__vss n1749__vss 25e-3
ri2242 n1666__vss n1750__vss 25e-3
ri2243 n1664__vss n1751__vss 500e-3
ri2244 n1706__vss n1713__vss 9.804e-3
ri2245 n1708__vss n1713__vss 8.333e-3
ri2246 n1710__vss n1713__vss 8.333e-3
ri2247 n1612__vss n1687__vss 125e-3
ri2248 n1637__vss n1687__vss 125e-3
ri2249 n1647__vss n1687__vss 125e-3
ri2250 n1600__vss n1687__vss 125e-3
ri2251 n1303__vss n1687__vss 125e-3
ri2252 n1559__vss n1687__vss 125e-3
ri2253 n1570__vss n1687__vss 125e-3
ri2254 n1656__vss n1687__vss 125e-3
ri2255 n1672__vss n1687__vss 125e-3
ri2256 n1669__vss n1687__vss 125e-3
ri2257 n1310__vss n1687__vss 125e-3
ri2258 n1681__vss n1687__vss 125e-3
ri2259 n1678__vss n1687__vss 125e-3
ri2260 n1886__vddio n1887__vddio 49.1e-3
ri2261 n1887__vddio n1888__vddio 2.546e-3
ri2262 n1888__vddio n1889__vddio 23.28e-3
ri2263 n1889__vddio n1890__vddio 26.19e-3
ri2264 n1890__vddio n1891__vddio 25.8e-3
ri2265 n1891__vddio n1892__vddio 24.53e-3
ri2266 n1892__vddio n1893__vddio 15.46e-3
ri2267 n1893__vddio n1894__vddio 15.28e-3
ri2268 n1894__vddio n1895__vddio 10.55e-3
ri2269 n1895__vddio n1896__vddio 24.73e-3
ri2270 n1896__vddio n1897__vddio 25.82e-3
ri2271 n1897__vddio n1898__vddio 10e-3
ri2272 n1898__vddio n1899__vddio 15.09e-3
ri2273 n1899__vddio n1900__vddio 15.64e-3
ri2274 n1900__vddio n1901__vddio 10.12e-3
ri2275 n1901__vddio n1902__vddio 24.71e-3
ri2276 n1902__vddio n1903__vddio 25.82e-3
ri2277 n1903__vddio n1904__vddio 10.37e-3
ri2278 n1904__vddio n1905__vddio 15.46e-3
ri2279 n1905__vddio n1906__vddio 15.28e-3
ri2280 n1906__vddio n1907__vddio 9.82e-3
ri2281 n1907__vddio n1908__vddio 25.46e-3
ri2282 n1908__vddio n1909__vddio 91.27e-3
ri2283 n1909__vddio n1910__vddio 115e-3
ri2284 n1910__vddio n1911__vddio 145.1e-3
ri2285 n1911__vddio n1912__vddio 12.09e-3
ri2286 n1912__vddio n1913__vddio 210.1e-3
ri2287 n1913__vddio n1914__vddio 12.09e-3
ri2288 n1914__vddio n1915__vddio 210.1e-3
ri2289 n1915__vddio n1916__vddio 12.09e-3
ri2290 n1916__vddio n1917__vddio 210.1e-3
ri2291 n1917__vddio n1918__vddio 12.09e-3
ri2292 n1918__vddio n1919__vddio 210.1e-3
ri2293 n1919__vddio n1920__vddio 12.09e-3
ri2294 n1920__vddio n1921__vddio 210.1e-3
ri2295 n1921__vddio n1922__vddio 12.09e-3
ri2296 n1922__vddio n1923__vddio 210.1e-3
ri2297 n1923__vddio n1924__vddio 12.09e-3
ri2298 n1924__vddio n1925__vddio 210.1e-3
ri2299 n1925__vddio n1926__vddio 12.09e-3
ri2300 n1926__vddio n1927__vddio 210.1e-3
ri2301 n1927__vddio n1928__vddio 12.09e-3
ri2302 n1928__vddio n1929__vddio 210.1e-3
ri2303 n1929__vddio n1930__vddio 12.09e-3
ri2304 n1930__vddio n1931__vddio 210.1e-3
ri2305 n1931__vddio n1932__vddio 12.09e-3
ri2306 n1932__vddio n1933__vddio 210.1e-3
ri2307 n1933__vddio n1934__vddio 12.09e-3
ri2308 n1934__vddio n1935__vddio 210.1e-3
ri2309 n1935__vddio n1936__vddio 12.09e-3
ri2310 n1936__vddio n1937__vddio 210.1e-3
ri2311 n1937__vddio n1938__vddio 12.09e-3
ri2312 n1938__vddio n1939__vddio 210.1e-3
ri2313 n1939__vddio n1940__vddio 12.09e-3
ri2314 n1940__vddio n1941__vddio 210.1e-3
ri2315 n1941__vddio n1595__vddio 57.95e-3
ri2316 n1813__vddio n1886__vddio 125e-3
ri2317 n1828__vddio n1888__vddio 125e-3
ri2318 n1879__vddio n1889__vddio 9.804e-3
ri2319 n1830__vddio n1890__vddio 125e-3
ri2320 n1792__vddio n1891__vddio 125e-3
ri2321 n1833__vddio n1893__vddio 125e-3
ri2322 n1881__vddio n1894__vddio 8.333e-3
ri2323 n1835__vddio n1895__vddio 125e-3
ri2324 n1837__vddio n1896__vddio 125e-3
ri2325 n1839__vddio n1897__vddio 125e-3
ri2326 n1841__vddio n1899__vddio 125e-3
ri2327 n1883__vddio n1900__vddio 8.333e-3
ri2328 n1843__vddio n1901__vddio 125e-3
ri2329 n1706__vddio n1902__vddio 125e-3
ri2330 n1846__vddio n1903__vddio 125e-3
ri2331 n1848__vddio n1905__vddio 125e-3
ri2332 n1885__vddio n1906__vddio 8.333e-3
ri2333 n1850__vddio n1907__vddio 125e-3
ri2334 n1852__vddio n1908__vddio 125e-3
ri2335 n1529__vddio n1910__vddio 16.67e-3
ri2336 n1533__vddio n1912__vddio 8.333e-3
ri2337 n1538__vddio n1914__vddio 8.333e-3
ri2338 n1543__vddio n1916__vddio 8.333e-3
ri2339 n1547__vddio n1918__vddio 8.333e-3
ri2340 n1551__vddio n1920__vddio 8.333e-3
ri2341 n1555__vddio n1922__vddio 8.333e-3
ri2342 n1559__vddio n1924__vddio 8.333e-3
ri2343 n1563__vddio n1926__vddio 8.333e-3
ri2344 n1567__vddio n1928__vddio 8.333e-3
ri2345 n1571__vddio n1930__vddio 8.333e-3
ri2346 n1575__vddio n1932__vddio 8.333e-3
ri2347 n1579__vddio n1934__vddio 8.333e-3
ri2348 n1583__vddio n1936__vddio 8.333e-3
ri2349 n1587__vddio n1938__vddio 8.333e-3
ri2350 n1591__vddio n1940__vddio 8.333e-3
ri2351 n78__i1__net3 n76__i1__net3 118.4e-3
ri2353 n76__i1__net3 n74__i1__net3 18.14e-3
ri2355 n74__i1__net3 n72__i1__net3 36.4e-3
ri2357 n72__i1__net3 n70__i1__net3 17.53e-3
ri2359 n70__i1__net3 n84__i1__net3 44.21e-3
ri2360 n84__i1__net3 n67__i1__net3 28.95e-3
ri2362 n84__i1__net3 n66__i1__net3 27.21e-3
rj1 n18__chipdriverout n26__chipdriverout 166.7e-3
rj2 n27__chipdriverout n19__chipdriverout 166.7e-3
rj3 n21__chipdriverout n28__chipdriverout 166.7e-3
rj4 n29__chipdriverout n22__chipdriverout 166.7e-3
rj5 n24__chipdriverout n30__chipdriverout 166.7e-3
rj6 n31__chipdriverout n14__chipdriverout 83.33e-3
rj7 n12__chipdriverout n32__chipdriverout 166.7e-3
rj8 n33__chipdriverout n11__chipdriverout 166.7e-3
rj9 n9__chipdriverout n34__chipdriverout 166.7e-3
rj10 n35__chipdriverout n8__chipdriverout 166.7e-3
rj11 n6__chipdriverout n36__chipdriverout 166.7e-3
rj12 n37__chipdriverout n5__chipdriverout 166.7e-3
rj13 n2__chipdriverout n38__chipdriverout 166.7e-3
rj14 n63__i1__i14__net1 n61__i1__i14__net1 125e-3
rj15 n63__i1__i14__net1 n62__i1__i14__net1 125e-3
rj16 n7__vss n10__vss 166.7e-3
rj17 n11__vss n6__vss 166.7e-3
rj18 n4__vss n12__vss 166.7e-3
rj19 n13__vss n3__vss 166.7e-3
rj20 n2__vddio n15__vddio 166.7e-3
rj21 n16__vddio n5__vddio 166.7e-3
rj22 n6__vddio n17__vddio 166.7e-3
rj23 n18__vddio n8__vddio 166.7e-3
rj24 n9__vddio n19__vddio 166.7e-3
rj25 n20__vddio n11__vddio 166.7e-3
rj26 n12__vddio n21__vddio 166.7e-3
rj27 n71__i1__i14__net1 n69__i1__i14__net1 125e-3
rj28 n70__i1__i14__net1 n71__i1__i14__net1 125e-3
rj29 n57__chipdriverout n65__chipdriverout 166.7e-3
rj30 n66__chipdriverout n58__chipdriverout 166.7e-3
rj31 n60__chipdriverout n67__chipdriverout 166.7e-3
rj32 n68__chipdriverout n61__chipdriverout 166.7e-3
rj33 n63__chipdriverout n69__chipdriverout 166.7e-3
rj34 n70__chipdriverout n40__chipdriverout 166.7e-3
rj35 n43__chipdriverout n71__chipdriverout 166.7e-3
rj36 n72__chipdriverout n44__chipdriverout 166.7e-3
rj37 n46__chipdriverout n73__chipdriverout 166.7e-3
rj38 n74__chipdriverout n47__chipdriverout 166.7e-3
rj39 n49__chipdriverout n75__chipdriverout 166.7e-3
rj40 n76__chipdriverout n50__chipdriverout 166.7e-3
rj41 n52__chipdriverout n77__chipdriverout 166.7e-3
rj42 n73__i1__i14__net1 n75__i1__i14__net1 125e-3
rj43 n75__i1__i14__net1 n74__i1__i14__net1 125e-3
rj44 n20__vss n23__vss 166.7e-3
rj45 n24__vss n19__vss 166.7e-3
rj46 n17__vss n25__vss 166.7e-3
rj47 n26__vss n16__vss 166.7e-3
rj48 n23__vddio n36__vddio 166.7e-3
rj49 n37__vddio n26__vddio 166.7e-3
rj50 n27__vddio n38__vddio 166.7e-3
rj51 n39__vddio n29__vddio 166.7e-3
rj52 n30__vddio n40__vddio 166.7e-3
rj53 n41__vddio n32__vddio 166.7e-3
rj54 n33__vddio n42__vddio 166.7e-3
rj55 n85__i1__i14__net1 n14__i1__i14__net1 250e-3
rj56 n16__i1__i14__net1 n85__i1__i14__net1 250e-3
rj57 n96__chipdriverout n104__chipdriverout 166.7e-3
rj58 n105__chipdriverout n97__chipdriverout 166.7e-3
rj59 n99__chipdriverout n106__chipdriverout 166.7e-3
rj60 n107__chipdriverout n100__chipdriverout 166.7e-3
rj61 n102__chipdriverout n108__chipdriverout 166.7e-3
rj62 n109__chipdriverout n79__chipdriverout 166.7e-3
rj63 n82__chipdriverout n110__chipdriverout 166.7e-3
rj64 n111__chipdriverout n83__chipdriverout 166.7e-3
rj65 n85__chipdriverout n112__chipdriverout 166.7e-3
rj66 n113__chipdriverout n86__chipdriverout 166.7e-3
rj67 n88__chipdriverout n114__chipdriverout 166.7e-3
rj68 n115__chipdriverout n89__chipdriverout 166.7e-3
rj69 n91__chipdriverout n116__chipdriverout 166.7e-3
rj70 n95__i1__i14__net1 n93__i1__i14__net1 125e-3
rj71 n94__i1__i14__net1 n95__i1__i14__net1 125e-3
rj72 n33__vss n36__vss 166.7e-3
rj73 n37__vss n32__vss 166.7e-3
rj74 n30__vss n38__vss 166.7e-3
rj75 n39__vss n29__vss 166.7e-3
rj76 n44__vddio n57__vddio 166.7e-3
rj77 n58__vddio n47__vddio 166.7e-3
rj78 n48__vddio n59__vddio 166.7e-3
rj79 n60__vddio n50__vddio 166.7e-3
rj80 n51__vddio n61__vddio 166.7e-3
rj81 n62__vddio n53__vddio 166.7e-3
rj82 n54__vddio n63__vddio 166.7e-3
rj84 n23__i5__clk4 n19__i5__clk4 383.3e-3
rj85 n19__i5__clk4 n22__i5__clk4 1.115
rj87 n103__i1__i14__net1 n101__i1__i14__net1 125e-3
rj88 n102__i1__i14__net1 n103__i1__i14__net1 125e-3
rj89 n135__chipdriverout n143__chipdriverout 166.7e-3
rj90 n144__chipdriverout n136__chipdriverout 166.7e-3
rj91 n138__chipdriverout n145__chipdriverout 166.7e-3
rj92 n146__chipdriverout n139__chipdriverout 166.7e-3
rj93 n141__chipdriverout n147__chipdriverout 166.7e-3
rj94 n148__chipdriverout n118__chipdriverout 166.7e-3
rj95 n121__chipdriverout n149__chipdriverout 166.7e-3
rj96 n150__chipdriverout n122__chipdriverout 166.7e-3
rj97 n124__chipdriverout n151__chipdriverout 166.7e-3
rj98 n152__chipdriverout n125__chipdriverout 166.7e-3
rj99 n127__chipdriverout n153__chipdriverout 166.7e-3
rj100 n154__chipdriverout n128__chipdriverout 166.7e-3
rj101 n130__chipdriverout n155__chipdriverout 166.7e-3
rj102 n10__i5__i7__i0__net1 n7__i5__i7__i0__net1 1
rj103 n7__i5__i7__i1__net1 n10__i5__i7__i1__net1 1
rj104 n109__i1__i14__net1 n111__i1__i14__net1 125e-3
rj105 n111__i1__i14__net1 n110__i1__i14__net1 125e-3
rj106 n46__vss n49__vss 166.7e-3
rj107 n50__vss n45__vss 166.7e-3
rj108 n43__vss n51__vss 166.7e-3
rj109 n52__vss n42__vss 166.7e-3
rj110 n69__vddio n82__vddio 166.7e-3
rj111 n83__vddio n72__vddio 166.7e-3
rj112 n73__vddio n84__vddio 166.7e-3
rj113 n85__vddio n75__vddio 166.7e-3
rj114 n76__vddio n86__vddio 166.7e-3
rj115 n87__vddio n78__vddio 166.7e-3
rj116 n79__vddio n88__vddio 166.7e-3
rj117 n7__x0 n6__x0 1.0037
rj118 n7__y0 n6__y0 1.0037
rj119 n119__i1__i14__net1 n117__i1__i14__net1 125e-3
rj120 n118__i1__i14__net1 n119__i1__i14__net1 125e-3
rj121 n182__chipdriverout n159__chipdriverout 166.7e-3
rj122 n160__chipdriverout n183__chipdriverout 166.7e-3
rj123 n184__chipdriverout n162__chipdriverout 166.7e-3
rj124 n163__chipdriverout n185__chipdriverout 166.7e-3
rj125 n186__chipdriverout n165__chipdriverout 166.7e-3
rj126 n168__chipdriverout n187__chipdriverout 166.7e-3
rj127 n188__chipdriverout n171__chipdriverout 166.7e-3
rj128 n172__chipdriverout n189__chipdriverout 166.7e-3
rj129 n190__chipdriverout n174__chipdriverout 166.7e-3
rj130 n175__chipdriverout n191__chipdriverout 166.7e-3
rj131 n192__chipdriverout n177__chipdriverout 166.7e-3
rj132 n178__chipdriverout n193__chipdriverout 166.7e-3
rj133 n194__chipdriverout n180__chipdriverout 166.7e-3
rj134 n121__i1__i14__net1 n34__i1__i14__net1 250e-3
rj135 n36__i1__i14__net1 n121__i1__i14__net1 250e-3
rj136 n62__vss n59__vss 166.7e-3
rj137 n58__vss n63__vss 166.7e-3
rj138 n64__vss n56__vss 166.7e-3
rj139 n55__vss n65__vss 166.7e-3
rj140 n109__vddio n96__vddio 166.7e-3
rj141 n99__vddio n110__vddio 166.7e-3
rj142 n111__vddio n100__vddio 166.7e-3
rj143 n102__vddio n112__vddio 166.7e-3
rj144 n113__vddio n103__vddio 166.7e-3
rj145 n105__vddio n114__vddio 166.7e-3
rj146 n115__vddio n106__vddio 166.7e-3
rj147 n129__i1__i14__net1 n135__i1__i14__net1 125e-3
rj148 n135__i1__i14__net1 n130__i1__i14__net1 125e-3
rj149 n221__chipdriverout n198__chipdriverout 166.7e-3
rj150 n199__chipdriverout n222__chipdriverout 166.7e-3
rj151 n223__chipdriverout n201__chipdriverout 166.7e-3
rj152 n202__chipdriverout n224__chipdriverout 166.7e-3
rj153 n225__chipdriverout n204__chipdriverout 166.7e-3
rj154 n207__chipdriverout n226__chipdriverout 166.7e-3
rj155 n227__chipdriverout n210__chipdriverout 166.7e-3
rj156 n211__chipdriverout n228__chipdriverout 166.7e-3
rj157 n229__chipdriverout n213__chipdriverout 166.7e-3
rj158 n214__chipdriverout n230__chipdriverout 166.7e-3
rj159 n231__chipdriverout n216__chipdriverout 166.7e-3
rj160 n217__chipdriverout n232__chipdriverout 166.7e-3
rj161 n233__chipdriverout n219__chipdriverout 166.7e-3
rj162 n139__i1__i14__net1 n137__i1__i14__net1 125e-3
rj163 n138__i1__i14__net1 n139__i1__i14__net1 125e-3
rj164 n75__vss n72__vss 166.7e-3
rj165 n71__vss n76__vss 166.7e-3
rj166 n77__vss n69__vss 166.7e-3
rj167 n68__vss n78__vss 166.7e-3
rj168 n130__vddio n117__vddio 166.7e-3
rj169 n120__vddio n131__vddio 166.7e-3
rj170 n132__vddio n121__vddio 166.7e-3
rj171 n123__vddio n133__vddio 166.7e-3
rj172 n134__vddio n124__vddio 166.7e-3
rj173 n126__vddio n135__vddio 166.7e-3
rj174 n136__vddio n127__vddio 166.7e-3
rj175 n149__i1__i14__net1 n151__i1__i14__net1 125e-3
rj176 n151__i1__i14__net1 n150__i1__i14__net1 125e-3
rj177 n260__chipdriverout n237__chipdriverout 166.7e-3
rj178 n238__chipdriverout n261__chipdriverout 166.7e-3
rj179 n262__chipdriverout n240__chipdriverout 166.7e-3
rj180 n241__chipdriverout n263__chipdriverout 166.7e-3
rj181 n264__chipdriverout n243__chipdriverout 166.7e-3
rj182 n246__chipdriverout n265__chipdriverout 166.7e-3
rj183 n266__chipdriverout n249__chipdriverout 166.7e-3
rj184 n250__chipdriverout n267__chipdriverout 166.7e-3
rj185 n268__chipdriverout n252__chipdriverout 166.7e-3
rj186 n253__chipdriverout n269__chipdriverout 166.7e-3
rj187 n270__chipdriverout n255__chipdriverout 166.7e-3
rj188 n256__chipdriverout n271__chipdriverout 166.7e-3
rj189 n272__chipdriverout n258__chipdriverout 166.7e-3
rj190 n32__i5__clk4 n30__i5__clk4 1.6189
rj192 n14__i5__i7__i0__net1 n13__i5__i7__i0__net1 1.5652
rj193 n13__i5__i7__i0__net1 n15__i5__i7__i0__net1 500e-3
rj194 n33__i5__clk4 n31__i5__clk4 1.6189
rj196 n14__i5__i7__i1__net1 n13__i5__i7__i1__net1 1.5652
rj197 n13__i5__i7__i1__net1 n15__i5__i7__i1__net1 500e-3
rj198 n153__i1__i14__net1 n155__i1__i14__net1 125e-3
rj199 n155__i1__i14__net1 n154__i1__i14__net1 125e-3
rj200 n88__vss n85__vss 166.7e-3
rj201 n84__vss n89__vss 166.7e-3
rj202 n90__vss n82__vss 166.7e-3
rj203 n81__vss n91__vss 166.7e-3
rj204 n151__vddio n138__vddio 166.7e-3
rj205 n141__vddio n152__vddio 166.7e-3
rj206 n153__vddio n142__vddio 166.7e-3
rj207 n144__vddio n154__vddio 166.7e-3
rj208 n155__vddio n145__vddio 166.7e-3
rj209 n147__vddio n156__vddio 166.7e-3
rj210 n157__vddio n148__vddio 166.7e-3
rj211 n165__i1__i14__net1 n167__i1__i14__net1 125e-3
rj212 n167__i1__i14__net1 n166__i1__i14__net1 125e-3
rj213 n10__reset n9__reset 573.1e-3
rj214 n11__reset n12__reset 1.0731
rj215 n299__chipdriverout n276__chipdriverout 166.7e-3
rj216 n277__chipdriverout n300__chipdriverout 166.7e-3
rj217 n301__chipdriverout n279__chipdriverout 166.7e-3
rj218 n280__chipdriverout n302__chipdriverout 166.7e-3
rj219 n303__chipdriverout n282__chipdriverout 166.7e-3
rj220 n285__chipdriverout n304__chipdriverout 166.7e-3
rj221 n305__chipdriverout n288__chipdriverout 166.7e-3
rj222 n289__chipdriverout n306__chipdriverout 166.7e-3
rj223 n307__chipdriverout n291__chipdriverout 166.7e-3
rj224 n292__chipdriverout n308__chipdriverout 166.7e-3
rj225 n309__chipdriverout n294__chipdriverout 166.7e-3
rj226 n295__chipdriverout n310__chipdriverout 166.7e-3
rj227 n311__chipdriverout n297__chipdriverout 166.7e-3
rj228 n58__i1__i14__net1 n170__i1__i14__net1 250e-3
rj229 n170__i1__i14__net1 n60__i1__i14__net1 250e-3
rj230 n6__i5__i7__x0out n2__i5__i7__x0out 1
rj231 n6__i5__i7__y0out n2__i5__i7__y0out 1
rj232 n98__vss n101__vss 166.7e-3
rj233 n102__vss n97__vss 166.7e-3
rj234 n95__vss n103__vss 166.7e-3
rj235 n104__vss n94__vss 166.7e-3
rj236 n159__vddio n172__vddio 166.7e-3
rj237 n173__vddio n162__vddio 166.7e-3
rj238 n163__vddio n174__vddio 166.7e-3
rj239 n175__vddio n165__vddio 166.7e-3
rj240 n166__vddio n176__vddio 166.7e-3
rj241 n177__vddio n168__vddio 166.7e-3
rj242 n169__vddio n178__vddio 166.7e-3
rj243 n183__i1__i14__net1 n181__i1__i14__net1 125e-3
rj244 n182__i1__i14__net1 n183__i1__i14__net1 125e-3
rj245 n5__x1 n6__x1 1.0019
rj246 n5__y1 n7__y1 1.0019
rj247 n315__chipdriverout n338__chipdriverout 166.7e-3
rj248 n339__chipdriverout n316__chipdriverout 166.7e-3
rj249 n318__chipdriverout n340__chipdriverout 166.7e-3
rj250 n341__chipdriverout n319__chipdriverout 166.7e-3
rj251 n321__chipdriverout n342__chipdriverout 166.7e-3
rj252 n343__chipdriverout n324__chipdriverout 166.7e-3
rj253 n327__chipdriverout n344__chipdriverout 166.7e-3
rj254 n345__chipdriverout n328__chipdriverout 166.7e-3
rj255 n330__chipdriverout n346__chipdriverout 166.7e-3
rj256 n347__chipdriverout n331__chipdriverout 166.7e-3
rj257 n333__chipdriverout n348__chipdriverout 166.7e-3
rj258 n349__chipdriverout n334__chipdriverout 166.7e-3
rj259 n336__chipdriverout n350__chipdriverout 166.7e-3
rj260 n189__i1__i14__net1 n191__i1__i14__net1 125e-3
rj261 n191__i1__i14__net1 n190__i1__i14__net1 125e-3
rj262 n111__vss n114__vss 166.7e-3
rj263 n115__vss n110__vss 166.7e-3
rj264 n108__vss n116__vss 166.7e-3
rj265 n117__vss n107__vss 166.7e-3
rj266 n180__vddio n193__vddio 166.7e-3
rj267 n194__vddio n183__vddio 166.7e-3
rj268 n184__vddio n195__vddio 166.7e-3
rj269 n196__vddio n186__vddio 166.7e-3
rj270 n187__vddio n197__vddio 166.7e-3
rj271 n198__vddio n189__vddio 166.7e-3
rj272 n190__vddio n199__vddio 166.7e-3
rj273 n193__i1__i14__net1 n82__i1__i14__net1 250e-3
rj274 n84__i1__i14__net1 n193__i1__i14__net1 250e-3
rj275 n354__chipdriverout n377__chipdriverout 166.7e-3
rj276 n378__chipdriverout n355__chipdriverout 166.7e-3
rj277 n357__chipdriverout n379__chipdriverout 166.7e-3
rj278 n380__chipdriverout n358__chipdriverout 166.7e-3
rj279 n360__chipdriverout n381__chipdriverout 166.7e-3
rj280 n382__chipdriverout n363__chipdriverout 166.7e-3
rj281 n366__chipdriverout n383__chipdriverout 166.7e-3
rj282 n384__chipdriverout n367__chipdriverout 166.7e-3
rj283 n369__chipdriverout n385__chipdriverout 166.7e-3
rj284 n386__chipdriverout n370__chipdriverout 166.7e-3
rj285 n372__chipdriverout n387__chipdriverout 166.7e-3
rj286 n388__chipdriverout n373__chipdriverout 166.7e-3
rj287 n375__chipdriverout n389__chipdriverout 166.7e-3
rj288 n90__i1__i14__net1 n206__i1__i14__net1 250e-3
rj289 n206__i1__i14__net1 n92__i1__i14__net1 250e-3
rj290 n124__vss n127__vss 166.7e-3
rj291 n128__vss n123__vss 166.7e-3
rj292 n121__vss n129__vss 166.7e-3
rj293 n130__vss n120__vss 166.7e-3
rj294 n211__vddio n224__vddio 166.7e-3
rj295 n225__vddio n214__vddio 166.7e-3
rj296 n215__vddio n226__vddio 166.7e-3
rj297 n227__vddio n217__vddio 166.7e-3
rj298 n218__vddio n228__vddio 166.7e-3
rj299 n229__vddio n220__vddio 166.7e-3
rj300 n221__vddio n230__vddio 166.7e-3
rj301 n215__i1__i14__net1 n213__i1__i14__net1 125e-3
rj302 n214__i1__i14__net1 n215__i1__i14__net1 125e-3
rj303 n393__chipdriverout n416__chipdriverout 166.7e-3
rj304 n417__chipdriverout n394__chipdriverout 166.7e-3
rj305 n396__chipdriverout n418__chipdriverout 166.7e-3
rj306 n419__chipdriverout n397__chipdriverout 166.7e-3
rj307 n399__chipdriverout n420__chipdriverout 166.7e-3
rj308 n421__chipdriverout n402__chipdriverout 166.7e-3
rj309 n405__chipdriverout n422__chipdriverout 166.7e-3
rj310 n423__chipdriverout n406__chipdriverout 166.7e-3
rj311 n408__chipdriverout n424__chipdriverout 166.7e-3
rj312 n425__chipdriverout n409__chipdriverout 166.7e-3
rj313 n411__chipdriverout n426__chipdriverout 166.7e-3
rj314 n427__chipdriverout n412__chipdriverout 166.7e-3
rj315 n414__chipdriverout n428__chipdriverout 166.7e-3
rj316 n223__i1__i14__net1 n221__i1__i14__net1 125e-3
rj317 n222__i1__i14__net1 n223__i1__i14__net1 125e-3
rj318 n50__i5__clk4 n44__i5__clk4 1.6189
rj320 n23__i5__i7__i0__net1 n20__i5__i7__i0__net1 2.0652
rj321 n20__i5__i7__i0__net1 n24__i5__i7__i0__net1 500e-3
rj322 n52__i5__clk4 n45__i5__clk4 1.6189
rj324 n23__i5__i7__i1__net1 n20__i5__i7__i1__net1 2.0652
rj325 n20__i5__i7__i1__net1 n24__i5__i7__i1__net1 500e-3
rj326 n131__vss n132__vss 166.7e-3
rj327 n133__vss n134__vss 166.7e-3
rj328 n135__vss n136__vss 166.7e-3
rj329 n137__vss n138__vss 166.7e-3
rj330 n231__vddio n232__vddio 166.7e-3
rj331 n233__vddio n234__vddio 166.7e-3
rj332 n235__vddio n236__vddio 166.7e-3
rj333 n237__vddio n238__vddio 166.7e-3
rj334 n239__vddio n240__vddio 166.7e-3
rj335 n241__vddio n242__vddio 166.7e-3
rj336 n243__vddio n244__vddio 166.7e-3
rj337 n231__i1__i14__net1 n229__i1__i14__net1 125e-3
rj338 n230__i1__i14__net1 n231__i1__i14__net1 125e-3
rj339 n432__chipdriverout n455__chipdriverout 166.7e-3
rj340 n456__chipdriverout n433__chipdriverout 166.7e-3
rj341 n435__chipdriverout n457__chipdriverout 166.7e-3
rj342 n458__chipdriverout n436__chipdriverout 166.7e-3
rj343 n438__chipdriverout n459__chipdriverout 166.7e-3
rj344 n460__chipdriverout n441__chipdriverout 166.7e-3
rj345 n444__chipdriverout n461__chipdriverout 166.7e-3
rj346 n462__chipdriverout n445__chipdriverout 166.7e-3
rj347 n447__chipdriverout n463__chipdriverout 166.7e-3
rj348 n464__chipdriverout n448__chipdriverout 166.7e-3
rj349 n450__chipdriverout n465__chipdriverout 166.7e-3
rj350 n466__chipdriverout n451__chipdriverout 166.7e-3
rj351 n453__chipdriverout n467__chipdriverout 166.7e-3
rj352 n22__reset n20__reset 573.1e-3
rj353 n23__reset n21__reset 573.1e-3
rj354 n233__i1__i14__net1 n235__i1__i14__net1 125e-3
rj355 n235__i1__i14__net1 n234__i1__i14__net1 125e-3
rj356 n150__vss n153__vss 166.7e-3
rj357 n154__vss n149__vss 166.7e-3
rj358 n147__vss n155__vss 166.7e-3
rj359 n156__vss n146__vss 166.7e-3
rj360 n253__vddio n266__vddio 166.7e-3
rj361 n267__vddio n256__vddio 166.7e-3
rj362 n257__vddio n268__vddio 166.7e-3
rj363 n269__vddio n259__vddio 166.7e-3
rj364 n260__vddio n270__vddio 166.7e-3
rj365 n271__vddio n262__vddio 166.7e-3
rj366 n263__vddio n272__vddio 166.7e-3
rj367 n2__i5__i7__x1out n6__i5__i7__x1out 1.0012
rj368 n247__i1__i14__net1 n245__i1__i14__net1 125e-3
rj369 n246__i1__i14__net1 n247__i1__i14__net1 125e-3
rj370 n2__i5__i7__y1out n6__i5__i7__y1out 1.0012
rj371 n486__chipdriverout n494__chipdriverout 166.7e-3
rj372 n495__chipdriverout n487__chipdriverout 166.7e-3
rj373 n489__chipdriverout n496__chipdriverout 166.7e-3
rj374 n497__chipdriverout n490__chipdriverout 166.7e-3
rj375 n492__chipdriverout n498__chipdriverout 166.7e-3
rj376 n499__chipdriverout n469__chipdriverout 166.7e-3
rj377 n472__chipdriverout n500__chipdriverout 166.7e-3
rj378 n501__chipdriverout n473__chipdriverout 166.7e-3
rj379 n475__chipdriverout n502__chipdriverout 166.7e-3
rj380 n503__chipdriverout n476__chipdriverout 166.7e-3
rj381 n478__chipdriverout n504__chipdriverout 166.7e-3
rj382 n505__chipdriverout n479__chipdriverout 166.7e-3
rj383 n481__chipdriverout n506__chipdriverout 166.7e-3
rj384 n7__x2 n6__x2 1.0027
rj385 n7__y2 n6__y2 1.0027
rj386 n142__i1__i14__net1 n250__i1__i14__net1 250e-3
rj387 n250__i1__i14__net1 n144__i1__i14__net1 250e-3
rj388 n166__vss n163__vss 166.7e-3
rj389 n162__vss n167__vss 166.7e-3
rj390 n168__vss n160__vss 166.7e-3
rj391 n159__vss n169__vss 166.7e-3
rj392 n297__vddio n284__vddio 166.7e-3
rj393 n287__vddio n298__vddio 166.7e-3
rj394 n299__vddio n288__vddio 166.7e-3
rj395 n290__vddio n300__vddio 166.7e-3
rj396 n301__vddio n291__vddio 166.7e-3
rj397 n293__vddio n302__vddio 166.7e-3
rj398 n303__vddio n294__vddio 166.7e-3
rj399 n263__i1__i14__net1 n261__i1__i14__net1 125e-3
rj400 n262__i1__i14__net1 n263__i1__i14__net1 125e-3
rj401 n507__chipdriverout n508__chipdriverout 166.7e-3
rj402 n509__chipdriverout n510__chipdriverout 166.7e-3
rj403 n511__chipdriverout n512__chipdriverout 166.7e-3
rj404 n513__chipdriverout n514__chipdriverout 166.7e-3
rj405 n515__chipdriverout n516__chipdriverout 166.7e-3
rj406 n517__chipdriverout n518__chipdriverout 166.7e-3
rj407 n519__chipdriverout n520__chipdriverout 166.7e-3
rj408 n521__chipdriverout n522__chipdriverout 166.7e-3
rj409 n523__chipdriverout n524__chipdriverout 166.7e-3
rj410 n525__chipdriverout n526__chipdriverout 166.7e-3
rj411 n527__chipdriverout n528__chipdriverout 166.7e-3
rj412 n529__chipdriverout n530__chipdriverout 166.7e-3
rj413 n531__chipdriverout n532__chipdriverout 166.7e-3
rj414 n265__i1__i14__net1 n267__i1__i14__net1 125e-3
rj415 n267__i1__i14__net1 n266__i1__i14__net1 125e-3
rj416 n170__vss n171__vss 166.7e-3
rj417 n172__vss n173__vss 166.7e-3
rj418 n174__vss n175__vss 166.7e-3
rj419 n176__vss n177__vss 166.7e-3
rj420 n304__vddio n305__vddio 166.7e-3
rj421 n306__vddio n307__vddio 166.7e-3
rj422 n308__vddio n309__vddio 166.7e-3
rj423 n310__vddio n311__vddio 166.7e-3
rj424 n312__vddio n313__vddio 166.7e-3
rj425 n314__vddio n315__vddio 166.7e-3
rj426 n316__vddio n317__vddio 166.7e-3
rj427 n277__i1__i14__net1 n162__i1__i14__net1 250e-3
rj428 n164__i1__i14__net1 n277__i1__i14__net1 250e-3
rj429 n546__chipdriverout n547__chipdriverout 166.7e-3
rj430 n548__chipdriverout n549__chipdriverout 166.7e-3
rj431 n550__chipdriverout n551__chipdriverout 166.7e-3
rj432 n552__chipdriverout n553__chipdriverout 166.7e-3
rj433 n554__chipdriverout n555__chipdriverout 166.7e-3
rj434 n556__chipdriverout n557__chipdriverout 166.7e-3
rj435 n558__chipdriverout n559__chipdriverout 166.7e-3
rj436 n560__chipdriverout n561__chipdriverout 166.7e-3
rj437 n562__chipdriverout n563__chipdriverout 166.7e-3
rj438 n564__chipdriverout n565__chipdriverout 166.7e-3
rj439 n566__chipdriverout n567__chipdriverout 166.7e-3
rj440 n568__chipdriverout n569__chipdriverout 166.7e-3
rj441 n570__chipdriverout n571__chipdriverout 166.7e-3
rj442 n283__i1__i14__net1 n281__i1__i14__net1 125e-3
rj443 n282__i1__i14__net1 n283__i1__i14__net1 125e-3
rj444 n189__vss n192__vss 166.7e-3
rj445 n193__vss n188__vss 166.7e-3
rj446 n186__vss n194__vss 166.7e-3
rj447 n195__vss n185__vss 166.7e-3
rj448 n326__vddio n339__vddio 166.7e-3
rj449 n340__vddio n329__vddio 166.7e-3
rj450 n330__vddio n341__vddio 166.7e-3
rj451 n342__vddio n332__vddio 166.7e-3
rj452 n333__vddio n343__vddio 166.7e-3
rj453 n344__vddio n335__vddio 166.7e-3
rj454 n336__vddio n345__vddio 166.7e-3
rj455 n60__i5__clk4 n58__i5__clk4 1.6189
rj457 n28__i5__i7__i0__net1 n27__i5__i7__i0__net1 1.5652
rj458 n27__i5__i7__i0__net1 n29__i5__i7__i0__net1 500e-3
rj459 n61__i5__clk4 n59__i5__clk4 1.6189
rj461 n28__i5__i7__i1__net1 n27__i5__i7__i1__net1 1.5652
rj462 n27__i5__i7__i1__net1 n29__i5__i7__i1__net1 500e-3
rj463 n289__i1__i14__net1 n291__i1__i14__net1 125e-3
rj464 n291__i1__i14__net1 n290__i1__i14__net1 125e-3
rj465 n603__chipdriverout n611__chipdriverout 166.7e-3
rj466 n612__chipdriverout n604__chipdriverout 166.7e-3
rj467 n606__chipdriverout n613__chipdriverout 166.7e-3
rj468 n614__chipdriverout n607__chipdriverout 166.7e-3
rj469 n609__chipdriverout n615__chipdriverout 166.7e-3
rj470 n616__chipdriverout n586__chipdriverout 166.7e-3
rj471 n589__chipdriverout n617__chipdriverout 166.7e-3
rj472 n618__chipdriverout n590__chipdriverout 166.7e-3
rj473 n592__chipdriverout n619__chipdriverout 166.7e-3
rj474 n620__chipdriverout n593__chipdriverout 166.7e-3
rj475 n595__chipdriverout n621__chipdriverout 166.7e-3
rj476 n622__chipdriverout n596__chipdriverout 166.7e-3
rj477 n598__chipdriverout n623__chipdriverout 166.7e-3
rj478 n186__i1__i14__net1 n298__i1__i14__net1 250e-3
rj479 n298__i1__i14__net1 n188__i1__i14__net1 250e-3
rj480 n28__reset n29__reset 1.0731
rj481 n30__reset n31__reset 1.0731
rj482 n196__vss n197__vss 166.7e-3
rj483 n198__vss n199__vss 166.7e-3
rj484 n200__vss n201__vss 166.7e-3
rj485 n202__vss n203__vss 166.7e-3
rj486 n346__vddio n347__vddio 166.7e-3
rj487 n348__vddio n349__vddio 166.7e-3
rj488 n350__vddio n351__vddio 166.7e-3
rj489 n352__vddio n353__vddio 166.7e-3
rj490 n354__vddio n355__vddio 166.7e-3
rj491 n356__vddio n357__vddio 166.7e-3
rj492 n358__vddio n359__vddio 166.7e-3
rj493 n309__i1__i14__net1 n311__i1__i14__net1 125e-3
rj494 n311__i1__i14__net1 n310__i1__i14__net1 125e-3
rj495 n9__i5__i7__x2out n5__i5__i7__x2out 1
rj496 n650__chipdriverout n642__chipdriverout 166.7e-3
rj497 n643__chipdriverout n651__chipdriverout 166.7e-3
rj498 n652__chipdriverout n645__chipdriverout 166.7e-3
rj499 n646__chipdriverout n653__chipdriverout 166.7e-3
rj500 n654__chipdriverout n648__chipdriverout 166.7e-3
rj501 n625__chipdriverout n655__chipdriverout 166.7e-3
rj502 n656__chipdriverout n628__chipdriverout 166.7e-3
rj503 n629__chipdriverout n657__chipdriverout 166.7e-3
rj504 n658__chipdriverout n631__chipdriverout 166.7e-3
rj505 n632__chipdriverout n659__chipdriverout 166.7e-3
rj506 n660__chipdriverout n634__chipdriverout 166.7e-3
rj507 n635__chipdriverout n661__chipdriverout 166.7e-3
rj508 n662__chipdriverout n637__chipdriverout 166.7e-3
rj509 n9__i5__i7__y2out n5__i5__i7__y2out 1
rj510 n202__i1__i14__net1 n318__i1__i14__net1 250e-3
rj511 n318__i1__i14__net1 n204__i1__i14__net1 250e-3
rj512 n5__x3 n6__x3 1.0027
rj513 n5__y3 n6__y3 1.0027
rj514 n209__vss n210__vss 166.7e-3
rj515 n211__vss n212__vss 166.7e-3
rj516 n213__vss n214__vss 166.7e-3
rj517 n215__vss n216__vss 166.7e-3
rj518 n367__vddio n368__vddio 166.7e-3
rj519 n369__vddio n370__vddio 166.7e-3
rj520 n371__vddio n372__vddio 166.7e-3
rj521 n373__vddio n374__vddio 166.7e-3
rj522 n375__vddio n376__vddio 166.7e-3
rj523 n377__vddio n378__vddio 166.7e-3
rj524 n379__vddio n380__vddio 166.7e-3
rj525 n321__i1__i14__net1 n323__i1__i14__net1 125e-3
rj526 n323__i1__i14__net1 n322__i1__i14__net1 125e-3
rj527 n689__chipdriverout n681__chipdriverout 166.7e-3
rj528 n682__chipdriverout n690__chipdriverout 166.7e-3
rj529 n691__chipdriverout n684__chipdriverout 166.7e-3
rj530 n685__chipdriverout n692__chipdriverout 166.7e-3
rj531 n693__chipdriverout n687__chipdriverout 166.7e-3
rj532 n664__chipdriverout n694__chipdriverout 166.7e-3
rj533 n695__chipdriverout n667__chipdriverout 166.7e-3
rj534 n668__chipdriverout n696__chipdriverout 166.7e-3
rj535 n697__chipdriverout n670__chipdriverout 166.7e-3
rj536 n671__chipdriverout n698__chipdriverout 166.7e-3
rj537 n699__chipdriverout n673__chipdriverout 166.7e-3
rj538 n674__chipdriverout n700__chipdriverout 166.7e-3
rj539 n701__chipdriverout n676__chipdriverout 166.7e-3
rj540 n331__i1__i14__net1 n329__i1__i14__net1 125e-3
rj541 n330__i1__i14__net1 n331__i1__i14__net1 125e-3
rj542 n222__vss n223__vss 166.7e-3
rj543 n224__vss n225__vss 166.7e-3
rj544 n226__vss n227__vss 166.7e-3
rj545 n228__vss n229__vss 166.7e-3
rj546 n388__vddio n389__vddio 166.7e-3
rj547 n390__vddio n391__vddio 166.7e-3
rj548 n392__vddio n393__vddio 166.7e-3
rj549 n394__vddio n395__vddio 166.7e-3
rj550 n396__vddio n397__vddio 166.7e-3
rj551 n398__vddio n399__vddio 166.7e-3
rj552 n400__vddio n401__vddio 166.7e-3
rj553 n337__i1__i14__net1 n339__i1__i14__net1 125e-3
rj554 n339__i1__i14__net1 n338__i1__i14__net1 125e-3
rj555 n728__chipdriverout n720__chipdriverout 166.7e-3
rj556 n721__chipdriverout n729__chipdriverout 166.7e-3
rj557 n730__chipdriverout n723__chipdriverout 166.7e-3
rj558 n724__chipdriverout n731__chipdriverout 166.7e-3
rj559 n732__chipdriverout n726__chipdriverout 166.7e-3
rj560 n703__chipdriverout n733__chipdriverout 166.7e-3
rj561 n734__chipdriverout n706__chipdriverout 166.7e-3
rj562 n707__chipdriverout n735__chipdriverout 166.7e-3
rj563 n736__chipdriverout n709__chipdriverout 166.7e-3
rj564 n710__chipdriverout n737__chipdriverout 166.7e-3
rj565 n738__chipdriverout n712__chipdriverout 166.7e-3
rj566 n713__chipdriverout n739__chipdriverout 166.7e-3
rj567 n740__chipdriverout n715__chipdriverout 166.7e-3
rj568 n349__i1__i14__net1 n351__i1__i14__net1 125e-3
rj569 n351__i1__i14__net1 n350__i1__i14__net1 125e-3
rj570 n235__vss n236__vss 166.7e-3
rj571 n237__vss n238__vss 166.7e-3
rj572 n239__vss n240__vss 166.7e-3
rj573 n241__vss n242__vss 166.7e-3
rj574 n409__vddio n410__vddio 166.7e-3
rj575 n411__vddio n412__vddio 166.7e-3
rj576 n413__vddio n414__vddio 166.7e-3
rj577 n415__vddio n416__vddio 166.7e-3
rj578 n417__vddio n418__vddio 166.7e-3
rj579 n419__vddio n420__vddio 166.7e-3
rj580 n421__vddio n422__vddio 166.7e-3
rj581 n355__i1__i14__net1 n353__i1__i14__net1 125e-3
rj582 n354__i1__i14__net1 n355__i1__i14__net1 125e-3
rj583 n74__i5__clk4 n64__i5__clk4 1.6189
rj585 n32__i5__i7__i0__net1 n30__i5__i7__i0__net1 1.5652
rj587 n75__i5__clk4 n68__i5__clk4 1.6189
rj589 n32__i5__i7__i1__net1 n30__i5__i7__i1__net1 1.5652
rj591 n759__chipdriverout n767__chipdriverout 166.7e-3
rj592 n768__chipdriverout n760__chipdriverout 166.7e-3
rj593 n762__chipdriverout n769__chipdriverout 166.7e-3
rj594 n770__chipdriverout n763__chipdriverout 166.7e-3
rj595 n765__chipdriverout n771__chipdriverout 166.7e-3
rj596 n772__chipdriverout n742__chipdriverout 166.7e-3
rj597 n745__chipdriverout n773__chipdriverout 166.7e-3
rj598 n774__chipdriverout n746__chipdriverout 166.7e-3
rj599 n748__chipdriverout n775__chipdriverout 166.7e-3
rj600 n776__chipdriverout n749__chipdriverout 166.7e-3
rj601 n751__chipdriverout n777__chipdriverout 166.7e-3
rj602 n778__chipdriverout n752__chipdriverout 166.7e-3
rj603 n754__chipdriverout n779__chipdriverout 166.7e-3
rj604 n367__i1__i14__net1 n365__i1__i14__net1 125e-3
rj605 n366__i1__i14__net1 n367__i1__i14__net1 125e-3
rj606 n248__vss n249__vss 166.7e-3
rj607 n250__vss n251__vss 166.7e-3
rj608 n252__vss n253__vss 166.7e-3
rj609 n254__vss n255__vss 166.7e-3
rj610 n434__vddio n435__vddio 166.7e-3
rj611 n436__vddio n437__vddio 166.7e-3
rj612 n438__vddio n439__vddio 166.7e-3
rj613 n440__vddio n441__vddio 166.7e-3
rj614 n442__vddio n443__vddio 166.7e-3
rj615 n444__vddio n445__vddio 166.7e-3
rj616 n446__vddio n447__vddio 166.7e-3
rj617 n33__reset n32__reset 573.1e-3
rj618 n34__reset n35__reset 1.0731
rj619 n369__i1__i14__net1 n371__i1__i14__net1 125e-3
rj620 n371__i1__i14__net1 n370__i1__i14__net1 125e-3
rj621 n806__chipdriverout n783__chipdriverout 166.7e-3
rj622 n784__chipdriverout n807__chipdriverout 166.7e-3
rj623 n808__chipdriverout n786__chipdriverout 166.7e-3
rj624 n787__chipdriverout n809__chipdriverout 166.7e-3
rj625 n810__chipdriverout n789__chipdriverout 166.7e-3
rj626 n792__chipdriverout n811__chipdriverout 166.7e-3
rj627 n812__chipdriverout n795__chipdriverout 166.7e-3
rj628 n796__chipdriverout n813__chipdriverout 166.7e-3
rj629 n814__chipdriverout n798__chipdriverout 166.7e-3
rj630 n799__chipdriverout n815__chipdriverout 166.7e-3
rj631 n816__chipdriverout n801__chipdriverout 166.7e-3
rj632 n802__chipdriverout n817__chipdriverout 166.7e-3
rj633 n818__chipdriverout n804__chipdriverout 166.7e-3
rj634 n383__i1__i14__net1 n377__i1__i14__net1 125e-3
rj635 n378__i1__i14__net1 n383__i1__i14__net1 125e-3
rj636 n9__i5__i7__x3out n5__i5__i7__x3out 1
rj637 n11__i5__i7__y3out n7__i5__i7__y3out 1
rj638 n267__vss n270__vss 166.7e-3
rj639 n271__vss n266__vss 166.7e-3
rj640 n264__vss n272__vss 166.7e-3
rj641 n273__vss n263__vss 166.7e-3
rj642 n462__vddio n475__vddio 166.7e-3
rj643 n476__vddio n465__vddio 166.7e-3
rj644 n466__vddio n477__vddio 166.7e-3
rj645 n478__vddio n468__vddio 166.7e-3
rj646 n469__vddio n479__vddio 166.7e-3
rj647 n480__vddio n471__vddio 166.7e-3
rj648 n472__vddio n481__vddio 166.7e-3
rj649 n387__i1__i14__net1 n385__i1__i14__net1 125e-3
rj650 n386__i1__i14__net1 n387__i1__i14__net1 125e-3
rj651 n845__chipdriverout n822__chipdriverout 166.7e-3
rj652 n823__chipdriverout n846__chipdriverout 166.7e-3
rj653 n847__chipdriverout n825__chipdriverout 166.7e-3
rj654 n826__chipdriverout n848__chipdriverout 166.7e-3
rj655 n849__chipdriverout n828__chipdriverout 166.7e-3
rj656 n831__chipdriverout n850__chipdriverout 166.7e-3
rj657 n851__chipdriverout n834__chipdriverout 166.7e-3
rj658 n835__chipdriverout n852__chipdriverout 166.7e-3
rj659 n853__chipdriverout n837__chipdriverout 166.7e-3
rj660 n838__chipdriverout n854__chipdriverout 166.7e-3
rj661 n855__chipdriverout n840__chipdriverout 166.7e-3
rj662 n841__chipdriverout n856__chipdriverout 166.7e-3
rj663 n857__chipdriverout n843__chipdriverout 166.7e-3
rj664 n286__i1__i14__net1 n398__i1__i14__net1 250e-3
rj665 n398__i1__i14__net1 n288__i1__i14__net1 250e-3
rj666 n280__vss n283__vss 166.7e-3
rj667 n284__vss n279__vss 166.7e-3
rj668 n277__vss n285__vss 166.7e-3
rj669 n286__vss n276__vss 166.7e-3
rj670 n483__vddio n496__vddio 166.7e-3
rj671 n497__vddio n486__vddio 166.7e-3
rj672 n487__vddio n498__vddio 166.7e-3
rj673 n499__vddio n489__vddio 166.7e-3
rj674 n490__vddio n500__vddio 166.7e-3
rj675 n501__vddio n492__vddio 166.7e-3
rj676 n493__vddio n502__vddio 166.7e-3
rj677 n403__i1__i14__net1 n401__i1__i14__net1 125e-3
rj678 n402__i1__i14__net1 n403__i1__i14__net1 125e-3
rj679 n16__i5__i7__y2out n14__i5__i7__y2out 565.9e-3
rj681 n16__i5__i7__y1out n13__i5__i7__y1out 565.5e-3
rj683 n873__chipdriverout n859__chipdriverout 166.7e-3
rj684 n862__chipdriverout n874__chipdriverout 166.7e-3
rj685 n875__chipdriverout n863__chipdriverout 166.7e-3
rj686 n865__chipdriverout n876__chipdriverout 166.7e-3
rj687 n877__chipdriverout n866__chipdriverout 166.7e-3
rj688 n868__chipdriverout n878__chipdriverout 166.7e-3
rj689 n879__chipdriverout n869__chipdriverout 166.7e-3
rj690 n871__chipdriverout n880__chipdriverout 166.7e-3
rj691 n11__i5__i7__x2out n13__i5__i7__x2out 404.1e-3
rj692 n12__i5__i7__x1out n13__i5__i7__x1out 433.4e-3
rj693 n884__chipdriverout n892__chipdriverout 166.7e-3
rj694 n893__chipdriverout n885__chipdriverout 166.7e-3
rj695 n887__chipdriverout n894__chipdriverout 166.7e-3
rj696 n895__chipdriverout n888__chipdriverout 166.7e-3
rj697 n890__chipdriverout n896__chipdriverout 166.7e-3
rj698 n411__i1__i14__net1 n409__i1__i14__net1 125e-3
rj699 n410__i1__i14__net1 n411__i1__i14__net1 125e-3
rj700 n517__vddio n504__vddio 166.7e-3
rj701 n507__vddio n518__vddio 166.7e-3
rj702 n519__vddio n508__vddio 166.7e-3
rj703 n510__vddio n520__vddio 166.7e-3
rj704 n521__vddio n511__vddio 166.7e-3
rj705 n513__vddio n522__vddio 166.7e-3
rj706 n523__vddio n514__vddio 166.7e-3
rj707 n287__vss n288__vss 166.7e-3
rj708 n289__vss n290__vss 166.7e-3
rj709 n298__vss n295__vss 166.7e-3
rj710 n294__vss n299__vss 166.7e-3
rj711 n9__i5__i7__xor2 n10__i5__i7__xor2 4.894e-3
rj712 n10__i5__i7__xor2 n8__i5__i7__xor2 160.4e-3
rj713 n6__i5__i7__xor2 n9__i5__i7__xor2 83.33e-3
rj714 n9__i5__i7__xor1 n10__i5__i7__xor1 4.894e-3
rj715 n10__i5__i7__xor1 n8__i5__i7__xor1 160.4e-3
rj716 n6__i5__i7__xor1 n9__i5__i7__xor1 83.33e-3
rj717 n417__i1__i14__net1 n419__i1__i14__net1 125e-3
rj718 n419__i1__i14__net1 n418__i1__i14__net1 125e-3
rj719 n923__chipdriverout n900__chipdriverout 166.7e-3
rj720 n901__chipdriverout n924__chipdriverout 166.7e-3
rj721 n925__chipdriverout n903__chipdriverout 166.7e-3
rj722 n904__chipdriverout n926__chipdriverout 166.7e-3
rj723 n927__chipdriverout n906__chipdriverout 166.7e-3
rj724 n909__chipdriverout n928__chipdriverout 166.7e-3
rj725 n929__chipdriverout n912__chipdriverout 166.7e-3
rj726 n913__chipdriverout n930__chipdriverout 166.7e-3
rj727 n931__chipdriverout n915__chipdriverout 166.7e-3
rj728 n916__chipdriverout n932__chipdriverout 166.7e-3
rj729 n933__chipdriverout n918__chipdriverout 166.7e-3
rj730 n919__chipdriverout n934__chipdriverout 166.7e-3
rj731 n935__chipdriverout n921__chipdriverout 166.7e-3
rj732 n429__i1__i14__net1 n314__i1__i14__net1 250e-3
rj733 n316__i1__i14__net1 n429__i1__i14__net1 250e-3
rj734 n300__vss n301__vss 166.7e-3
rj735 n302__vss n303__vss 166.7e-3
rj736 n304__vss n305__vss 166.7e-3
rj737 n306__vss n307__vss 166.7e-3
rj738 n538__vddio n525__vddio 166.7e-3
rj739 n528__vddio n539__vddio 166.7e-3
rj740 n540__vddio n529__vddio 166.7e-3
rj741 n531__vddio n541__vddio 166.7e-3
rj742 n542__vddio n532__vddio 166.7e-3
rj743 n534__vddio n543__vddio 166.7e-3
rj744 n544__vddio n535__vddio 166.7e-3
rj745 n437__i1__i14__net1 n439__i1__i14__net1 125e-3
rj746 n439__i1__i14__net1 n438__i1__i14__net1 125e-3
rj747 n962__chipdriverout n939__chipdriverout 166.7e-3
rj748 n940__chipdriverout n963__chipdriverout 166.7e-3
rj749 n964__chipdriverout n942__chipdriverout 166.7e-3
rj750 n943__chipdriverout n965__chipdriverout 166.7e-3
rj751 n966__chipdriverout n945__chipdriverout 166.7e-3
rj752 n948__chipdriverout n967__chipdriverout 166.7e-3
rj753 n968__chipdriverout n951__chipdriverout 166.7e-3
rj754 n952__chipdriverout n969__chipdriverout 166.7e-3
rj755 n970__chipdriverout n954__chipdriverout 166.7e-3
rj756 n955__chipdriverout n971__chipdriverout 166.7e-3
rj757 n972__chipdriverout n957__chipdriverout 166.7e-3
rj758 n958__chipdriverout n973__chipdriverout 166.7e-3
rj759 n974__chipdriverout n960__chipdriverout 166.7e-3
rj760 n445__i1__i14__net1 n334__i1__i14__net1 250e-3
rj761 n336__i1__i14__net1 n445__i1__i14__net1 250e-3
rj762 n313__vss n314__vss 166.7e-3
rj763 n315__vss n316__vss 166.7e-3
rj764 n317__vss n318__vss 166.7e-3
rj765 n319__vss n320__vss 166.7e-3
rj766 n545__vddio n546__vddio 166.7e-3
rj767 n547__vddio n548__vddio 166.7e-3
rj768 n549__vddio n550__vddio 166.7e-3
rj769 n551__vddio n552__vddio 166.7e-3
rj770 n553__vddio n554__vddio 166.7e-3
rj771 n555__vddio n556__vddio 166.7e-3
rj772 n557__vddio n558__vddio 166.7e-3
rj773 n453__i1__i14__net1 n455__i1__i14__net1 125e-3
rj774 n455__i1__i14__net1 n454__i1__i14__net1 125e-3
rj775 n975__chipdriverout n976__chipdriverout 166.7e-3
rj776 n977__chipdriverout n978__chipdriverout 166.7e-3
rj777 n979__chipdriverout n980__chipdriverout 166.7e-3
rj778 n981__chipdriverout n982__chipdriverout 166.7e-3
rj779 n983__chipdriverout n984__chipdriverout 166.7e-3
rj780 n985__chipdriverout n986__chipdriverout 166.7e-3
rj781 n987__chipdriverout n988__chipdriverout 166.7e-3
rj782 n989__chipdriverout n990__chipdriverout 166.7e-3
rj783 n991__chipdriverout n992__chipdriverout 166.7e-3
rj784 n993__chipdriverout n994__chipdriverout 166.7e-3
rj785 n995__chipdriverout n996__chipdriverout 166.7e-3
rj786 n997__chipdriverout n998__chipdriverout 166.7e-3
rj787 n999__chipdriverout n1000__chipdriverout 166.7e-3
rj788 n463__i1__i14__net1 n461__i1__i14__net1 125e-3
rj789 n462__i1__i14__net1 n463__i1__i14__net1 125e-3
rj790 n326__vss n327__vss 166.7e-3
rj791 n328__vss n329__vss 166.7e-3
rj792 n330__vss n331__vss 166.7e-3
rj793 n332__vss n333__vss 166.7e-3
rj794 n590__vddio n577__vddio 166.7e-3
rj795 n580__vddio n591__vddio 166.7e-3
rj796 n592__vddio n581__vddio 166.7e-3
rj797 n583__vddio n593__vddio 166.7e-3
rj798 n594__vddio n584__vddio 166.7e-3
rj799 n586__vddio n595__vddio 166.7e-3
rj800 n596__vddio n587__vddio 166.7e-3
rj801 n14__i5__i7__y3out n13__i5__i7__y3out 390e-3
rj802 n13__i5__i7__y3out n12__i5__i7__y3out 175.9e-3
rj803 n16__i5__i7__y0out n13__i5__i7__y0out 565.5e-3
rj805 n11__i5__i7__x3out n13__i5__i7__x3out 421.2e-3
rj806 n12__i5__i7__x0out n13__i5__i7__x0out 423.6e-3
rj807 n469__i1__i14__net1 n357__i1__i14__net1 250e-3
rj808 n359__i1__i14__net1 n469__i1__i14__net1 250e-3
rj809 n1040__chipdriverout n1017__chipdriverout 166.7e-3
rj810 n1018__chipdriverout n1041__chipdriverout 166.7e-3
rj811 n1042__chipdriverout n1020__chipdriverout 166.7e-3
rj812 n1021__chipdriverout n1043__chipdriverout 166.7e-3
rj813 n1044__chipdriverout n1023__chipdriverout 166.7e-3
rj814 n1026__chipdriverout n1045__chipdriverout 166.7e-3
rj815 n1046__chipdriverout n1029__chipdriverout 166.7e-3
rj816 n1030__chipdriverout n1047__chipdriverout 166.7e-3
rj817 n1048__chipdriverout n1032__chipdriverout 166.7e-3
rj818 n1033__chipdriverout n1049__chipdriverout 166.7e-3
rj819 n1050__chipdriverout n1035__chipdriverout 166.7e-3
rj820 n1036__chipdriverout n1051__chipdriverout 166.7e-3
rj821 n1052__chipdriverout n1038__chipdriverout 166.7e-3
rj822 n475__i1__i14__net1 n473__i1__i14__net1 125e-3
rj823 n474__i1__i14__net1 n475__i1__i14__net1 125e-3
rj824 n339__vss n340__vss 166.7e-3
rj825 n341__vss n342__vss 166.7e-3
rj826 n343__vss n344__vss 166.7e-3
rj827 n345__vss n346__vss 166.7e-3
rj828 n597__vddio n598__vddio 166.7e-3
rj829 n599__vddio n600__vddio 166.7e-3
rj830 n601__vddio n602__vddio 166.7e-3
rj831 n603__vddio n604__vddio 166.7e-3
rj832 n605__vddio n606__vddio 166.7e-3
rj833 n607__vddio n608__vddio 166.7e-3
rj834 n609__vddio n610__vddio 166.7e-3
rj835 n485__i1__i14__net1 n487__i1__i14__net1 125e-3
rj836 n487__i1__i14__net1 n486__i1__i14__net1 125e-3
rj837 n1079__chipdriverout n1056__chipdriverout 166.7e-3
rj838 n1057__chipdriverout n1080__chipdriverout 166.7e-3
rj839 n1081__chipdriverout n1059__chipdriverout 166.7e-3
rj840 n1060__chipdriverout n1082__chipdriverout 166.7e-3
rj841 n1083__chipdriverout n1062__chipdriverout 166.7e-3
rj842 n1065__chipdriverout n1084__chipdriverout 166.7e-3
rj843 n1085__chipdriverout n1068__chipdriverout 166.7e-3
rj844 n1069__chipdriverout n1086__chipdriverout 166.7e-3
rj845 n1087__chipdriverout n1071__chipdriverout 166.7e-3
rj846 n1072__chipdriverout n1088__chipdriverout 166.7e-3
rj847 n1089__chipdriverout n1074__chipdriverout 166.7e-3
rj848 n1075__chipdriverout n1090__chipdriverout 166.7e-3
rj849 n1091__chipdriverout n1077__chipdriverout 166.7e-3
rj850 n491__i1__i14__net1 n489__i1__i14__net1 125e-3
rj851 n490__i1__i14__net1 n491__i1__i14__net1 125e-3
rj852 n361__vss n358__vss 166.7e-3
rj853 n357__vss n362__vss 166.7e-3
rj854 n363__vss n355__vss 166.7e-3
rj855 n354__vss n364__vss 166.7e-3
rj856 n632__vddio n619__vddio 166.7e-3
rj857 n622__vddio n633__vddio 166.7e-3
rj858 n634__vddio n623__vddio 166.7e-3
rj859 n625__vddio n635__vddio 166.7e-3
rj860 n636__vddio n626__vddio 166.7e-3
rj861 n628__vddio n637__vddio 166.7e-3
rj862 n638__vddio n629__vddio 166.7e-3
rj863 n501__i1__i14__net1 n503__i1__i14__net1 125e-3
rj864 n503__i1__i14__net1 n502__i1__i14__net1 125e-3
rj865 n1092__chipdriverout n1093__chipdriverout 166.7e-3
rj866 n1094__chipdriverout n1095__chipdriverout 166.7e-3
rj867 n1096__chipdriverout n1097__chipdriverout 166.7e-3
rj868 n1098__chipdriverout n1099__chipdriverout 166.7e-3
rj869 n1100__chipdriverout n1101__chipdriverout 166.7e-3
rj870 n1102__chipdriverout n1103__chipdriverout 166.7e-3
rj871 n1104__chipdriverout n1105__chipdriverout 166.7e-3
rj872 n1106__chipdriverout n1107__chipdriverout 166.7e-3
rj873 n1108__chipdriverout n1109__chipdriverout 166.7e-3
rj874 n1110__chipdriverout n1111__chipdriverout 166.7e-3
rj875 n1112__chipdriverout n1113__chipdriverout 166.7e-3
rj876 n1114__chipdriverout n1115__chipdriverout 166.7e-3
rj877 n1116__chipdriverout n1117__chipdriverout 166.7e-3
rj878 n17__i5__i7__xor2 n15__i5__i7__xor2 500e-3
rj879 n15__i5__i7__xor1 n17__i5__i7__xor1 500e-3
rj880 n511__i1__i14__net1 n509__i1__i14__net1 125e-3
rj881 n510__i1__i14__net1 n511__i1__i14__net1 125e-3
rj882 n365__vss n366__vss 166.7e-3
rj883 n367__vss n368__vss 166.7e-3
rj884 n369__vss n370__vss 166.7e-3
rj885 n371__vss n372__vss 166.7e-3
rj886 n663__vddio n650__vddio 166.7e-3
rj887 n653__vddio n664__vddio 166.7e-3
rj888 n665__vddio n654__vddio 166.7e-3
rj889 n656__vddio n666__vddio 166.7e-3
rj890 n667__vddio n657__vddio 166.7e-3
rj891 n659__vddio n668__vddio 166.7e-3
rj892 n669__vddio n660__vddio 166.7e-3
rj893 n517__i1__i14__net1 n519__i1__i14__net1 125e-3
rj894 n519__i1__i14__net1 n518__i1__i14__net1 125e-3
rj895 n1157__chipdriverout n1134__chipdriverout 166.7e-3
rj896 n1135__chipdriverout n1158__chipdriverout 166.7e-3
rj897 n1159__chipdriverout n1137__chipdriverout 166.7e-3
rj898 n1138__chipdriverout n1160__chipdriverout 166.7e-3
rj899 n1161__chipdriverout n1140__chipdriverout 166.7e-3
rj900 n1143__chipdriverout n1162__chipdriverout 166.7e-3
rj901 n1163__chipdriverout n1146__chipdriverout 166.7e-3
rj902 n1147__chipdriverout n1164__chipdriverout 166.7e-3
rj903 n1165__chipdriverout n1149__chipdriverout 166.7e-3
rj904 n1150__chipdriverout n1166__chipdriverout 166.7e-3
rj905 n1167__chipdriverout n1152__chipdriverout 166.7e-3
rj906 n1153__chipdriverout n1168__chipdriverout 166.7e-3
rj907 n1169__chipdriverout n1155__chipdriverout 166.7e-3
rj908 n521__i1__i14__net1 n414__i1__i14__net1 250e-3
rj909 n416__i1__i14__net1 n521__i1__i14__net1 250e-3
rj910 n378__vss n379__vss 166.7e-3
rj911 n380__vss n381__vss 166.7e-3
rj912 n382__vss n383__vss 166.7e-3
rj913 n384__vss n385__vss 166.7e-3
rj914 n670__vddio n671__vddio 166.7e-3
rj915 n672__vddio n673__vddio 166.7e-3
rj916 n674__vddio n675__vddio 166.7e-3
rj917 n676__vddio n677__vddio 166.7e-3
rj918 n678__vddio n679__vddio 166.7e-3
rj919 n680__vddio n681__vddio 166.7e-3
rj920 n682__vddio n683__vddio 166.7e-3
rj921 n11__i5__i7__i5__net1 n10__i5__i7__i5__net1 125e-3
rj922 n10__i5__i7__i4__net1 n11__i5__i7__i4__net1 125e-3
rj923 n535__i1__i14__net1 n533__i1__i14__net1 125e-3
rj924 n534__i1__i14__net1 n535__i1__i14__net1 125e-3
rj925 n1196__chipdriverout n1173__chipdriverout 166.7e-3
rj926 n1174__chipdriverout n1197__chipdriverout 166.7e-3
rj927 n1198__chipdriverout n1176__chipdriverout 166.7e-3
rj928 n1177__chipdriverout n1199__chipdriverout 166.7e-3
rj929 n1200__chipdriverout n1179__chipdriverout 166.7e-3
rj930 n1182__chipdriverout n1201__chipdriverout 166.7e-3
rj931 n1202__chipdriverout n1185__chipdriverout 166.7e-3
rj932 n1186__chipdriverout n1203__chipdriverout 166.7e-3
rj933 n1204__chipdriverout n1188__chipdriverout 166.7e-3
rj934 n1189__chipdriverout n1205__chipdriverout 166.7e-3
rj935 n1206__chipdriverout n1191__chipdriverout 166.7e-3
rj936 n1192__chipdriverout n1207__chipdriverout 166.7e-3
rj937 n1208__chipdriverout n1194__chipdriverout 166.7e-3
rj938 n6__i5__i7__net47 n7__i5__i7__net47 250e-3
rj939 n4__i5__i7__net44 n5__i5__i7__net44 250e-3
rj940 n539__i1__i14__net1 n537__i1__i14__net1 125e-3
rj941 n538__i1__i14__net1 n539__i1__i14__net1 125e-3
rj942 n400__vss n397__vss 166.7e-3
rj943 n396__vss n401__vss 166.7e-3
rj944 n402__vss n394__vss 166.7e-3
rj945 n393__vss n403__vss 166.7e-3
rj946 n705__vddio n692__vddio 166.7e-3
rj947 n695__vddio n706__vddio 166.7e-3
rj948 n707__vddio n696__vddio 166.7e-3
rj949 n698__vddio n708__vddio 166.7e-3
rj950 n709__vddio n699__vddio 166.7e-3
rj951 n701__vddio n710__vddio 166.7e-3
rj952 n711__vddio n702__vddio 166.7e-3
rj953 n18__i5__i7__xor2 n19__i5__i7__xor2 250e-3
rj954 n18__i5__i7__xor1 n19__i5__i7__xor1 250e-3
rj955 n549__i1__i14__net1 n551__i1__i14__net1 125e-3
rj956 n551__i1__i14__net1 n550__i1__i14__net1 125e-3
rj957 n1212__chipdriverout n1235__chipdriverout 166.7e-3
rj958 n1236__chipdriverout n1213__chipdriverout 166.7e-3
rj959 n1215__chipdriverout n1237__chipdriverout 166.7e-3
rj960 n1238__chipdriverout n1216__chipdriverout 166.7e-3
rj961 n1218__chipdriverout n1239__chipdriverout 166.7e-3
rj962 n1240__chipdriverout n1221__chipdriverout 166.7e-3
rj963 n1224__chipdriverout n1241__chipdriverout 166.7e-3
rj964 n1242__chipdriverout n1225__chipdriverout 166.7e-3
rj965 n1227__chipdriverout n1243__chipdriverout 166.7e-3
rj966 n1244__chipdriverout n1228__chipdriverout 166.7e-3
rj967 n1230__chipdriverout n1245__chipdriverout 166.7e-3
rj968 n1246__chipdriverout n1231__chipdriverout 166.7e-3
rj969 n1233__chipdriverout n1247__chipdriverout 166.7e-3
rj970 n557__i1__i14__net1 n559__i1__i14__net1 125e-3
rj971 n559__i1__i14__net1 n558__i1__i14__net1 125e-3
rj972 n17__i5__i7__xor3 n18__i5__i7__xor3 246.1e-3
rj973 n18__i5__i7__xor3 n19__i5__i7__xor3 308.7e-3
rj974 n19__i5__i7__xor3 n20__i5__i7__xor3 434.2e-3
rj975 n19__i5__i7__xor3 n21__i5__i7__xor3 126.5e-3
rj977 n20__i5__i7__xor3 n6__i5__i7__xor3 165.3e-3
rj978 n21__i5__i7__xor3 n9__i5__i7__xor3 206.8e-3
rj979 n15__i5__i7__xor3 n18__i5__i7__xor3 125e-3
rj980 n8__i5__i7__xor3 n20__i5__i7__xor3 83.33e-3
rj981 n17__i5__i7__xor0 n18__i5__i7__xor0 246.1e-3
rj982 n18__i5__i7__xor0 n19__i5__i7__xor0 308.7e-3
rj983 n19__i5__i7__xor0 n20__i5__i7__xor0 434.2e-3
rj984 n19__i5__i7__xor0 n21__i5__i7__xor0 126.5e-3
rj986 n20__i5__i7__xor0 n6__i5__i7__xor0 165.3e-3
rj987 n21__i5__i7__xor0 n9__i5__i7__xor0 206.8e-3
rj988 n15__i5__i7__xor0 n18__i5__i7__xor0 125e-3
rj989 n8__i5__i7__xor0 n20__i5__i7__xor0 83.33e-3
rj990 n413__vss n410__vss 166.7e-3
rj991 n409__vss n414__vss 166.7e-3
rj992 n415__vss n407__vss 166.7e-3
rj993 n406__vss n416__vss 166.7e-3
rj994 n726__vddio n713__vddio 166.7e-3
rj995 n716__vddio n727__vddio 166.7e-3
rj996 n728__vddio n717__vddio 166.7e-3
rj997 n719__vddio n729__vddio 166.7e-3
rj998 n730__vddio n720__vddio 166.7e-3
rj999 n722__vddio n731__vddio 166.7e-3
rj1000 n732__vddio n723__vddio 166.7e-3
rj1001 n565__i1__i14__net1 n567__i1__i14__net1 125e-3
rj1002 n567__i1__i14__net1 n566__i1__i14__net1 125e-3
rj1003 n1274__chipdriverout n1251__chipdriverout 166.7e-3
rj1004 n1252__chipdriverout n1275__chipdriverout 166.7e-3
rj1005 n1276__chipdriverout n1254__chipdriverout 166.7e-3
rj1006 n1255__chipdriverout n1277__chipdriverout 166.7e-3
rj1007 n1278__chipdriverout n1257__chipdriverout 166.7e-3
rj1008 n1260__chipdriverout n1279__chipdriverout 166.7e-3
rj1009 n1280__chipdriverout n1263__chipdriverout 166.7e-3
rj1010 n1264__chipdriverout n1281__chipdriverout 166.7e-3
rj1011 n1282__chipdriverout n1266__chipdriverout 166.7e-3
rj1012 n1267__chipdriverout n1283__chipdriverout 166.7e-3
rj1013 n1284__chipdriverout n1269__chipdriverout 166.7e-3
rj1014 n1270__chipdriverout n1285__chipdriverout 166.7e-3
rj1015 n1286__chipdriverout n1272__chipdriverout 166.7e-3
rj1016 n573__i1__i14__net1 n575__i1__i14__net1 125e-3
rj1017 n575__i1__i14__net1 n574__i1__i14__net1 125e-3
rj1018 n14__i5__i7__i5__net1 n12__i5__i7__i5__net1 500e-3
rj1019 n12__i5__i7__i4__net1 n14__i5__i7__i4__net1 500e-3
rj1020 n423__vss n426__vss 166.7e-3
rj1021 n427__vss n422__vss 166.7e-3
rj1022 n420__vss n428__vss 166.7e-3
rj1023 n429__vss n419__vss 166.7e-3
rj1024 n734__vddio n747__vddio 166.7e-3
rj1025 n748__vddio n737__vddio 166.7e-3
rj1026 n738__vddio n749__vddio 166.7e-3
rj1027 n750__vddio n740__vddio 166.7e-3
rj1028 n741__vddio n751__vddio 166.7e-3
rj1029 n752__vddio n743__vddio 166.7e-3
rj1030 n744__vddio n753__vddio 166.7e-3
rj1032 n13__i5__i7__net51 n10__i5__i7__net51 157.3e-3
rj1033 n12__i5__i7__net51 n13__i5__i7__net51 83.33e-3
rj1034 n583__i1__i14__net1 n581__i1__i14__net1 125e-3
rj1035 n582__i1__i14__net1 n583__i1__i14__net1 125e-3
rj1036 n1290__chipdriverout n1313__chipdriverout 166.7e-3
rj1037 n1314__chipdriverout n1291__chipdriverout 166.7e-3
rj1038 n1293__chipdriverout n1315__chipdriverout 166.7e-3
rj1039 n1316__chipdriverout n1294__chipdriverout 166.7e-3
rj1040 n1296__chipdriverout n1317__chipdriverout 166.7e-3
rj1041 n1318__chipdriverout n1299__chipdriverout 166.7e-3
rj1042 n1302__chipdriverout n1319__chipdriverout 166.7e-3
rj1043 n1320__chipdriverout n1303__chipdriverout 166.7e-3
rj1044 n1305__chipdriverout n1321__chipdriverout 166.7e-3
rj1045 n1322__chipdriverout n1306__chipdriverout 166.7e-3
rj1046 n1308__chipdriverout n1323__chipdriverout 166.7e-3
rj1047 n1324__chipdriverout n1309__chipdriverout 166.7e-3
rj1048 n1311__chipdriverout n1325__chipdriverout 166.7e-3
rj1049 n478__i1__i14__net1 n586__i1__i14__net1 250e-3
rj1050 n586__i1__i14__net1 n480__i1__i14__net1 250e-3
rj1051 n430__vss n431__vss 166.7e-3
rj1052 n432__vss n433__vss 166.7e-3
rj1053 n434__vss n435__vss 166.7e-3
rj1054 n436__vss n437__vss 166.7e-3
rj1055 n755__vddio n768__vddio 166.7e-3
rj1056 n769__vddio n758__vddio 166.7e-3
rj1057 n759__vddio n770__vddio 166.7e-3
rj1058 n771__vddio n761__vddio 166.7e-3
rj1059 n762__vddio n772__vddio 166.7e-3
rj1060 n773__vddio n764__vddio 166.7e-3
rj1061 n765__vddio n774__vddio 166.7e-3
rj1062 n599__i1__i14__net1 n597__i1__i14__net1 125e-3
rj1063 n598__i1__i14__net1 n599__i1__i14__net1 125e-3
rj1064 n15__i5__i7__net51 n17__i5__i7__net51 500e-3
rj1065 n1352__chipdriverout n1329__chipdriverout 166.7e-3
rj1066 n1330__chipdriverout n1353__chipdriverout 166.7e-3
rj1067 n1354__chipdriverout n1332__chipdriverout 166.7e-3
rj1068 n1333__chipdriverout n1355__chipdriverout 166.7e-3
rj1069 n1356__chipdriverout n1335__chipdriverout 166.7e-3
rj1070 n1338__chipdriverout n1357__chipdriverout 166.7e-3
rj1071 n1358__chipdriverout n1341__chipdriverout 166.7e-3
rj1072 n1342__chipdriverout n1359__chipdriverout 166.7e-3
rj1073 n1360__chipdriverout n1344__chipdriverout 166.7e-3
rj1074 n1345__chipdriverout n1361__chipdriverout 166.7e-3
rj1075 n1362__chipdriverout n1347__chipdriverout 166.7e-3
rj1076 n1348__chipdriverout n1363__chipdriverout 166.7e-3
rj1077 n1364__chipdriverout n1350__chipdriverout 166.7e-3
rj1078 n601__i1__i14__net1 n603__i1__i14__net1 125e-3
rj1079 n603__i1__i14__net1 n602__i1__i14__net1 125e-3
rj1080 n449__vss n452__vss 166.7e-3
rj1081 n453__vss n448__vss 166.7e-3
rj1082 n446__vss n454__vss 166.7e-3
rj1083 n455__vss n445__vss 166.7e-3
rj1084 n776__vddio n789__vddio 166.7e-3
rj1085 n790__vddio n779__vddio 166.7e-3
rj1086 n780__vddio n791__vddio 166.7e-3
rj1087 n792__vddio n782__vddio 166.7e-3
rj1088 n783__vddio n793__vddio 166.7e-3
rj1089 n794__vddio n785__vddio 166.7e-3
rj1090 n786__vddio n795__vddio 166.7e-3
rj1091 n615__i1__i14__net1 n613__i1__i14__net1 125e-3
rj1092 n614__i1__i14__net1 n615__i1__i14__net1 125e-3
rj1093 n12__i5__i7__net47 n11__i5__i7__net47 494e-3
rj1094 n11__i5__i7__net47 n10__i5__i7__net47 71.92e-3
rj1095 n1368__chipdriverout n1391__chipdriverout 166.7e-3
rj1096 n1392__chipdriverout n1369__chipdriverout 166.7e-3
rj1097 n1371__chipdriverout n1393__chipdriverout 166.7e-3
rj1098 n1394__chipdriverout n1372__chipdriverout 166.7e-3
rj1099 n1374__chipdriverout n1395__chipdriverout 166.7e-3
rj1100 n1396__chipdriverout n1377__chipdriverout 166.7e-3
rj1101 n1380__chipdriverout n1397__chipdriverout 166.7e-3
rj1102 n1398__chipdriverout n1381__chipdriverout 166.7e-3
rj1103 n1383__chipdriverout n1399__chipdriverout 166.7e-3
rj1104 n1400__chipdriverout n1384__chipdriverout 166.7e-3
rj1105 n1386__chipdriverout n1401__chipdriverout 166.7e-3
rj1106 n1402__chipdriverout n1387__chipdriverout 166.7e-3
rj1107 n1389__chipdriverout n1403__chipdriverout 166.7e-3
rj1108 n8__i5__i7__net44 n9__i5__i7__net44 779.6e-3
rj1109 n623__i1__i14__net1 n621__i1__i14__net1 125e-3
rj1110 n622__i1__i14__net1 n623__i1__i14__net1 125e-3
rj1111 n3__i5__i7__i6__net1 n8__i5__i7__i6__net1 250e-3
rj1112 n462__vss n465__vss 166.7e-3
rj1113 n466__vss n461__vss 166.7e-3
rj1114 n459__vss n467__vss 166.7e-3
rj1115 n468__vss n458__vss 166.7e-3
rj1116 n801__vddio n814__vddio 166.7e-3
rj1117 n815__vddio n804__vddio 166.7e-3
rj1118 n805__vddio n816__vddio 166.7e-3
rj1119 n817__vddio n807__vddio 166.7e-3
rj1120 n808__vddio n818__vddio 166.7e-3
rj1121 n819__vddio n810__vddio 166.7e-3
rj1122 n811__vddio n820__vddio 166.7e-3
rj1123 n627__i1__i14__net1 n625__i1__i14__net1 125e-3
rj1124 n626__i1__i14__net1 n627__i1__i14__net1 125e-3
rj1125 n4__i5__i7__net46 n5__i5__i7__net46 250e-3
rj1126 n1430__chipdriverout n1407__chipdriverout 166.7e-3
rj1127 n1408__chipdriverout n1431__chipdriverout 166.7e-3
rj1128 n1432__chipdriverout n1410__chipdriverout 166.7e-3
rj1129 n1411__chipdriverout n1433__chipdriverout 166.7e-3
rj1130 n1434__chipdriverout n1413__chipdriverout 166.7e-3
rj1131 n1416__chipdriverout n1435__chipdriverout 166.7e-3
rj1132 n1436__chipdriverout n1419__chipdriverout 166.7e-3
rj1133 n1420__chipdriverout n1437__chipdriverout 166.7e-3
rj1134 n1438__chipdriverout n1422__chipdriverout 166.7e-3
rj1135 n1423__chipdriverout n1439__chipdriverout 166.7e-3
rj1136 n1440__chipdriverout n1425__chipdriverout 166.7e-3
rj1137 n1426__chipdriverout n1441__chipdriverout 166.7e-3
rj1138 n1442__chipdriverout n1428__chipdriverout 166.7e-3
rj1139 n635__i1__i14__net1 n633__i1__i14__net1 125e-3
rj1140 n634__i1__i14__net1 n635__i1__i14__net1 125e-3
rj1141 n18__i5__i7__net44 n12__i5__i7__net44 1
rj1142 n18__i5__i7__net51 n19__i5__i7__net51 250e-3
rj1143 n469__vss n470__vss 166.7e-3
rj1144 n471__vss n472__vss 166.7e-3
rj1145 n473__vss n474__vss 166.7e-3
rj1146 n475__vss n476__vss 166.7e-3
rj1147 n827__vddio n828__vddio 166.7e-3
rj1148 n829__vddio n830__vddio 166.7e-3
rj1149 n831__vddio n832__vddio 166.7e-3
rj1150 n833__vddio n834__vddio 166.7e-3
rj1151 n835__vddio n836__vddio 166.7e-3
rj1152 n837__vddio n838__vddio 166.7e-3
rj1153 n839__vddio n840__vddio 166.7e-3
rj1154 n530__i1__i14__net1 n642__i1__i14__net1 250e-3
rj1155 n642__i1__i14__net1 n532__i1__i14__net1 250e-3
rj1156 n17__i5__i7__net50 n18__i5__i7__net50 246.1e-3
rj1157 n18__i5__i7__net50 n19__i5__i7__net50 438.9e-3
rj1158 n19__i5__i7__net50 n20__i5__i7__net50 409.5e-3
rj1159 n20__i5__i7__net50 n8__i5__i7__net50 165.3e-3
rj1160 n19__i5__i7__net50 n9__i5__i7__net50 208.8e-3
rj1161 n15__i5__i7__net50 n18__i5__i7__net50 125e-3
rj1162 n6__i5__i7__net50 n20__i5__i7__net50 83.33e-3
rj1163 n1445__chipdriverout n1446__chipdriverout 166.7e-3
rj1164 n1447__chipdriverout n1448__chipdriverout 166.7e-3
rj1165 n1449__chipdriverout n1450__chipdriverout 166.7e-3
rj1166 n1451__chipdriverout n1452__chipdriverout 166.7e-3
rj1167 n1453__chipdriverout n1454__chipdriverout 166.7e-3
rj1168 n1455__chipdriverout n1456__chipdriverout 166.7e-3
rj1169 n1457__chipdriverout n1458__chipdriverout 166.7e-3
rj1170 n1459__chipdriverout n1460__chipdriverout 166.7e-3
rj1171 n1461__chipdriverout n1462__chipdriverout 166.7e-3
rj1172 n1463__chipdriverout n1464__chipdriverout 166.7e-3
rj1173 n1465__chipdriverout n1466__chipdriverout 166.7e-3
rj1174 n1467__chipdriverout n1468__chipdriverout 166.7e-3
rj1175 n1469__chipdriverout n1470__chipdriverout 166.7e-3
rj1176 n655__i1__i14__net1 n653__i1__i14__net1 125e-3
rj1177 n654__i1__i14__net1 n655__i1__i14__net1 125e-3
rj1178 n491__vss n488__vss 166.7e-3
rj1179 n487__vss n492__vss 166.7e-3
rj1180 n493__vss n485__vss 166.7e-3
rj1181 n484__vss n494__vss 166.7e-3
rj1182 n862__vddio n849__vddio 166.7e-3
rj1183 n852__vddio n863__vddio 166.7e-3
rj1184 n864__vddio n853__vddio 166.7e-3
rj1185 n855__vddio n865__vddio 166.7e-3
rj1186 n866__vddio n856__vddio 166.7e-3
rj1187 n858__vddio n867__vddio 166.7e-3
rj1188 n868__vddio n859__vddio 166.7e-3
rj1189 n663__i1__i14__net1 n661__i1__i14__net1 125e-3
rj1190 n662__i1__i14__net1 n663__i1__i14__net1 125e-3
rj1191 n1501__chipdriverout n1524__chipdriverout 166.7e-3
rj1192 n1525__chipdriverout n1502__chipdriverout 166.7e-3
rj1193 n1504__chipdriverout n1526__chipdriverout 166.7e-3
rj1194 n1527__chipdriverout n1505__chipdriverout 166.7e-3
rj1195 n1507__chipdriverout n1528__chipdriverout 166.7e-3
rj1196 n1529__chipdriverout n1510__chipdriverout 166.7e-3
rj1197 n1513__chipdriverout n1530__chipdriverout 166.7e-3
rj1198 n1531__chipdriverout n1514__chipdriverout 166.7e-3
rj1199 n1516__chipdriverout n1532__chipdriverout 166.7e-3
rj1200 n1533__chipdriverout n1517__chipdriverout 166.7e-3
rj1201 n1519__chipdriverout n1534__chipdriverout 166.7e-3
rj1202 n1535__chipdriverout n1520__chipdriverout 166.7e-3
rj1203 n1522__chipdriverout n1536__chipdriverout 166.7e-3
rj1204 n14__i5__i7__i6__net1 n12__i5__i7__i6__net1 500e-3
rj1205 n665__i1__i14__net1 n554__i1__i14__net1 250e-3
rj1206 n556__i1__i14__net1 n665__i1__i14__net1 250e-3
rj1207 n8__i5__r0 n10__i5__r0 161.5e-3
rj1208 n10__i5__r0 n9__i5__r0 2.416e-3
rj1209 n6__i5__r0 n10__i5__r0 83.33e-3
rj1210 n495__vss n496__vss 166.7e-3
rj1211 n497__vss n498__vss 166.7e-3
rj1212 n499__vss n500__vss 166.7e-3
rj1213 n501__vss n502__vss 166.7e-3
rj1214 n869__vddio n870__vddio 166.7e-3
rj1215 n871__vddio n872__vddio 166.7e-3
rj1216 n873__vddio n874__vddio 166.7e-3
rj1217 n875__vddio n876__vddio 166.7e-3
rj1218 n877__vddio n878__vddio 166.7e-3
rj1219 n879__vddio n880__vddio 166.7e-3
rj1220 n881__vddio n882__vddio 166.7e-3
rj1221 n12__i5__i7__net46 n13__i5__i7__net46 910.2e-3
rj1222 n677__i1__i14__net1 n562__i1__i14__net1 250e-3
rj1223 n564__i1__i14__net1 n677__i1__i14__net1 250e-3
rj1224 n16__i5__clk_buf n17__i5__clk_buf 500e-3
rj1225 n1541__chipdriverout n1564__chipdriverout 166.7e-3
rj1226 n1565__chipdriverout n1542__chipdriverout 166.7e-3
rj1227 n1544__chipdriverout n1566__chipdriverout 166.7e-3
rj1228 n1567__chipdriverout n1545__chipdriverout 166.7e-3
rj1229 n1547__chipdriverout n1568__chipdriverout 166.7e-3
rj1230 n1569__chipdriverout n1550__chipdriverout 166.7e-3
rj1231 n1553__chipdriverout n1570__chipdriverout 166.7e-3
rj1232 n1571__chipdriverout n1554__chipdriverout 166.7e-3
rj1233 n1556__chipdriverout n1572__chipdriverout 166.7e-3
rj1234 n1573__chipdriverout n1557__chipdriverout 166.7e-3
rj1235 n1559__chipdriverout n1574__chipdriverout 166.7e-3
rj1236 n1575__chipdriverout n1560__chipdriverout 166.7e-3
rj1237 n1562__chipdriverout n1576__chipdriverout 166.7e-3
rj1238 n681__i1__i14__net1 n570__i1__i14__net1 250e-3
rj1239 n572__i1__i14__net1 n681__i1__i14__net1 250e-3
rj1240 n6__i5__r1 n5__i5__r1 117.6e-3
rj1241 n6__i5__r1 n3__i5__r1 131e-3
rj1242 n514__vss n517__vss 166.7e-3
rj1243 n518__vss n513__vss 166.7e-3
rj1244 n511__vss n519__vss 166.7e-3
rj1245 n520__vss n510__vss 166.7e-3
rj1246 n891__vddio n914__vddio 166.7e-3
rj1247 n915__vddio n894__vddio 166.7e-3
rj1248 n895__vddio n916__vddio 166.7e-3
rj1249 n917__vddio n897__vddio 166.7e-3
rj1250 n898__vddio n918__vddio 166.7e-3
rj1251 n919__vddio n900__vddio 166.7e-3
rj1252 n901__vddio n920__vddio 166.7e-3
rj1253 n695__i1__i14__net1 n693__i1__i14__net1 125e-3
rj1254 n694__i1__i14__net1 n695__i1__i14__net1 125e-3
rj1255 n1581__chipdriverout n1604__chipdriverout 166.7e-3
rj1256 n1605__chipdriverout n1582__chipdriverout 166.7e-3
rj1257 n1584__chipdriverout n1606__chipdriverout 166.7e-3
rj1258 n1607__chipdriverout n1585__chipdriverout 166.7e-3
rj1259 n1587__chipdriverout n1608__chipdriverout 166.7e-3
rj1260 n1609__chipdriverout n1590__chipdriverout 166.7e-3
rj1261 n1593__chipdriverout n1610__chipdriverout 166.7e-3
rj1262 n1611__chipdriverout n1594__chipdriverout 166.7e-3
rj1263 n1596__chipdriverout n1612__chipdriverout 166.7e-3
rj1264 n1613__chipdriverout n1597__chipdriverout 166.7e-3
rj1265 n1599__chipdriverout n1614__chipdriverout 166.7e-3
rj1266 n1615__chipdriverout n1600__chipdriverout 166.7e-3
rj1267 n1602__chipdriverout n1616__chipdriverout 166.7e-3
rj1268 n15__i5__i6__net31 n12__i5__i6__net31 500e-3
rj1269 n590__i1__i14__net1 n698__i1__i14__net1 250e-3
rj1270 n698__i1__i14__net1 n592__i1__i14__net1 250e-3
rj1271 n530__vss n527__vss 166.7e-3
rj1272 n526__vss n531__vss 166.7e-3
rj1273 n532__vss n524__vss 166.7e-3
rj1274 n523__vss n533__vss 166.7e-3
rj1275 n935__vddio n922__vddio 166.7e-3
rj1276 n925__vddio n936__vddio 166.7e-3
rj1277 n937__vddio n926__vddio 166.7e-3
rj1278 n928__vddio n938__vddio 166.7e-3
rj1279 n939__vddio n929__vddio 166.7e-3
rj1280 n931__vddio n940__vddio 166.7e-3
rj1281 n941__vddio n932__vddio 166.7e-3
rj1282 n709__i1__i14__net1 n711__i1__i14__net1 125e-3
rj1283 n711__i1__i14__net1 n710__i1__i14__net1 125e-3
rj1284 n21__i5__i7__i7__net1 n22__i5__i7__i7__net1 940.4e-3
rj1285 n22__i5__i7__i7__net1 n23__i5__i7__i7__net1 628.1e-3
rj1286 n23__i5__i7__i7__net1 n24__i5__i7__i7__net1 292.2e-3
rj1287 n24__i5__i7__i7__net1 n16__i5__i7__i7__net1 22.04e-3
rj1288 n24__i5__i7__i7__net1 n25__i5__i7__i7__net1 693.5e-3
rj1289 n25__i5__i7__i7__net1 n13__i5__i7__i7__net1 106.4e-3
rj1290 n25__i5__i7__i7__net1 n11__i5__i7__i7__net1 141.9e-3
rj1291 n19__i5__i7__i7__net1 n23__i5__i7__i7__net1 250e-3
rj1292 n1635__chipdriverout n1643__chipdriverout 166.7e-3
rj1293 n1644__chipdriverout n1636__chipdriverout 166.7e-3
rj1294 n1638__chipdriverout n1645__chipdriverout 166.7e-3
rj1295 n1646__chipdriverout n1639__chipdriverout 166.7e-3
rj1296 n1641__chipdriverout n1647__chipdriverout 166.7e-3
rj1297 n1648__chipdriverout n1618__chipdriverout 166.7e-3
rj1298 n1621__chipdriverout n1649__chipdriverout 166.7e-3
rj1299 n1650__chipdriverout n1622__chipdriverout 166.7e-3
rj1300 n1624__chipdriverout n1651__chipdriverout 166.7e-3
rj1301 n1652__chipdriverout n1625__chipdriverout 166.7e-3
rj1302 n1627__chipdriverout n1653__chipdriverout 166.7e-3
rj1303 n1654__chipdriverout n1628__chipdriverout 166.7e-3
rj1304 n1630__chipdriverout n1655__chipdriverout 166.7e-3
rj1305 n719__i1__i14__net1 n717__i1__i14__net1 125e-3
rj1306 n718__i1__i14__net1 n719__i1__i14__net1 125e-3
rj1307 n44__vdd n46__vdd 1.2455
rj1308 n540__vss n543__vss 166.7e-3
rj1309 n544__vss n539__vss 166.7e-3
rj1310 n537__vss n545__vss 166.7e-3
rj1311 n546__vss n536__vss 166.7e-3
rj1312 n943__vddio n956__vddio 166.7e-3
rj1313 n957__vddio n946__vddio 166.7e-3
rj1314 n947__vddio n958__vddio 166.7e-3
rj1315 n959__vddio n949__vddio 166.7e-3
rj1316 n950__vddio n960__vddio 166.7e-3
rj1317 n961__vddio n952__vddio 166.7e-3
rj1318 n953__vddio n962__vddio 166.7e-3
rj1319 n15__shift n16__shift 1.0669
rj1320 n16__shift n13__shift 28.1e-3
rj1321 n9__shift n16__shift 500e-3
rj1323 n47__vdd n49__vdd 440.7e-3
rj1325 n49__vdd n51__vdd 440.7e-3
rj1327 n51__vdd n53__vdd 440.7e-3
rj1329 n53__vdd n55__vdd 440.7e-3
rj1331 n55__vdd n57__vdd 440.7e-3
rj1333 n57__vdd n59__vdd 440.7e-3
rj1335 n59__vdd n61__vdd 440.7e-3
rj1337 n61__vdd n63__vdd 440.7e-3
rj1339 n63__vdd n65__vdd 440.7e-3
rj1340 n65__vdd n66__vdd 12.5e-3
rj1341 n723__i1__i14__net1 n721__i1__i14__net1 125e-3
rj1342 n722__i1__i14__net1 n723__i1__i14__net1 125e-3
rj1343 n1674__chipdriverout n1682__chipdriverout 166.7e-3
rj1344 n1683__chipdriverout n1675__chipdriverout 166.7e-3
rj1345 n1677__chipdriverout n1684__chipdriverout 166.7e-3
rj1346 n1685__chipdriverout n1678__chipdriverout 166.7e-3
rj1347 n1680__chipdriverout n1686__chipdriverout 166.7e-3
rj1348 n1687__chipdriverout n1657__chipdriverout 166.7e-3
rj1349 n1660__chipdriverout n1688__chipdriverout 166.7e-3
rj1350 n1689__chipdriverout n1661__chipdriverout 166.7e-3
rj1351 n1663__chipdriverout n1690__chipdriverout 166.7e-3
rj1352 n1691__chipdriverout n1664__chipdriverout 166.7e-3
rj1353 n1666__chipdriverout n1692__chipdriverout 166.7e-3
rj1354 n1693__chipdriverout n1667__chipdriverout 166.7e-3
rj1355 n1669__chipdriverout n1694__chipdriverout 166.7e-3
rj1356 n725__i1__i14__net1 n727__i1__i14__net1 125e-3
rj1357 n727__i1__i14__net1 n726__i1__i14__net1 125e-3
rj1358 n4__i5__r2 n6__i5__r2 333.3e-3
rj1359 n562__vss n559__vss 166.7e-3
rj1360 n558__vss n563__vss 166.7e-3
rj1361 n564__vss n556__vss 166.7e-3
rj1362 n555__vss n565__vss 166.7e-3
rj1363 n977__vddio n964__vddio 166.7e-3
rj1364 n967__vddio n978__vddio 166.7e-3
rj1365 n979__vddio n968__vddio 166.7e-3
rj1366 n970__vddio n980__vddio 166.7e-3
rj1367 n981__vddio n971__vddio 166.7e-3
rj1368 n973__vddio n982__vddio 166.7e-3
rj1369 n983__vddio n974__vddio 166.7e-3
rj1370 n731__i1__i14__net1 n729__i1__i14__net1 125e-3
rj1371 n730__i1__i14__net1 n731__i1__i14__net1 125e-3
rj1372 n1721__chipdriverout n1713__chipdriverout 166.7e-3
rj1373 n1714__chipdriverout n1722__chipdriverout 166.7e-3
rj1374 n1723__chipdriverout n1716__chipdriverout 166.7e-3
rj1375 n1717__chipdriverout n1724__chipdriverout 166.7e-3
rj1376 n1725__chipdriverout n1719__chipdriverout 166.7e-3
rj1377 n1696__chipdriverout n1726__chipdriverout 166.7e-3
rj1378 n1727__chipdriverout n1699__chipdriverout 166.7e-3
rj1379 n1700__chipdriverout n1728__chipdriverout 166.7e-3
rj1380 n1729__chipdriverout n1702__chipdriverout 166.7e-3
rj1381 n1703__chipdriverout n1730__chipdriverout 166.7e-3
rj1382 n1731__chipdriverout n1705__chipdriverout 166.7e-3
rj1383 n1706__chipdriverout n1732__chipdriverout 166.7e-3
rj1384 n1733__chipdriverout n1708__chipdriverout 166.7e-3
rj1385 n15__i5__i6__net30 n9__i5__i6__net30 588.1e-3
rj1386 n735__i1__i14__net1 n733__i1__i14__net1 125e-3
rj1387 n734__i1__i14__net1 n735__i1__i14__net1 125e-3
rj1388 n572__vss n575__vss 166.7e-3
rj1389 n576__vss n571__vss 166.7e-3
rj1390 n569__vss n577__vss 166.7e-3
rj1391 n578__vss n568__vss 166.7e-3
rj1392 n985__vddio n998__vddio 166.7e-3
rj1393 n999__vddio n988__vddio 166.7e-3
rj1394 n989__vddio n1000__vddio 166.7e-3
rj1395 n1001__vddio n991__vddio 166.7e-3
rj1396 n992__vddio n1002__vddio 166.7e-3
rj1397 n1003__vddio n994__vddio 166.7e-3
rj1398 n995__vddio n1004__vddio 166.7e-3
rj1399 n739__i1__i14__net1 n737__i1__i14__net1 125e-3
rj1400 n738__i1__i14__net1 n739__i1__i14__net1 125e-3
rj1401 n27__i5__clk_buf n12__i5__clk_buf 1
rj1402 n1752__chipdriverout n1760__chipdriverout 166.7e-3
rj1403 n1761__chipdriverout n1753__chipdriverout 166.7e-3
rj1404 n1755__chipdriverout n1762__chipdriverout 166.7e-3
rj1405 n1763__chipdriverout n1756__chipdriverout 166.7e-3
rj1406 n1758__chipdriverout n1764__chipdriverout 166.7e-3
rj1407 n1765__chipdriverout n1735__chipdriverout 166.7e-3
rj1408 n1738__chipdriverout n1766__chipdriverout 166.7e-3
rj1409 n1767__chipdriverout n1739__chipdriverout 166.7e-3
rj1410 n1741__chipdriverout n1768__chipdriverout 166.7e-3
rj1411 n1769__chipdriverout n1742__chipdriverout 166.7e-3
rj1412 n1744__chipdriverout n1770__chipdriverout 166.7e-3
rj1413 n1771__chipdriverout n1745__chipdriverout 166.7e-3
rj1414 n1747__chipdriverout n1772__chipdriverout 166.7e-3
rj1415 n23__i5__i7__net46 n19__i5__i7__net46 198.7e-3
rj1416 n19__i5__i7__net46 n18__i5__i7__net46 98.66e-3
rj1417 n741__i1__i14__net1 n743__i1__i14__net1 125e-3
rj1418 n743__i1__i14__net1 n742__i1__i14__net1 125e-3
rj1419 n9__i5__i6__i2__net25 n6__i5__i6__i2__net25 176.5e-3
rj1420 n6__i5__i6__i2__net25 n3__i5__i6__i2__net25 178.9e-3
rj1421 n6__i5__i6__i2__net21 n9__i5__i6__i2__net21 494e-3
rj1422 n9__i5__i6__i2__net21 n2__i5__i6__i2__net21 236.9e-3
rj1423 n9__i5__i6__i2__net21 n3__i5__i6__i2__net21 278.9e-3
rj1424 n27__i5__i7__i7__net1 n28__i5__i7__i7__net1 1
rj1425 n579__vss n580__vss 166.7e-3
rj1426 n581__vss n582__vss 166.7e-3
rj1427 n583__vss n584__vss 166.7e-3
rj1428 n585__vss n586__vss 166.7e-3
rj1429 n1005__vddio n1006__vddio 166.7e-3
rj1430 n1007__vddio n1008__vddio 166.7e-3
rj1431 n1009__vddio n1010__vddio 166.7e-3
rj1432 n1011__vddio n1012__vddio 166.7e-3
rj1433 n1013__vddio n1014__vddio 166.7e-3
rj1434 n1015__vddio n1016__vddio 166.7e-3
rj1435 n1017__vddio n1018__vddio 166.7e-3
rj1436 n19__i5__i7__net44 n22__i5__i7__net44 718.6e-3
rj1437 n22__i5__i7__net44 n21__i5__i7__net44 218.8e-3
rj1438 n745__i1__i14__net1 n747__i1__i14__net1 125e-3
rj1439 n747__i1__i14__net1 n746__i1__i14__net1 125e-3
rj1440 n1799__chipdriverout n1791__chipdriverout 166.7e-3
rj1441 n1792__chipdriverout n1800__chipdriverout 166.7e-3
rj1442 n1801__chipdriverout n1794__chipdriverout 166.7e-3
rj1443 n1795__chipdriverout n1802__chipdriverout 166.7e-3
rj1444 n1803__chipdriverout n1797__chipdriverout 166.7e-3
rj1445 n1774__chipdriverout n1804__chipdriverout 166.7e-3
rj1446 n1805__chipdriverout n1777__chipdriverout 166.7e-3
rj1447 n1778__chipdriverout n1806__chipdriverout 166.7e-3
rj1448 n1807__chipdriverout n1780__chipdriverout 166.7e-3
rj1449 n1781__chipdriverout n1808__chipdriverout 166.7e-3
rj1450 n1809__chipdriverout n1783__chipdriverout 166.7e-3
rj1451 n1784__chipdriverout n1810__chipdriverout 166.7e-3
rj1452 n1811__chipdriverout n1786__chipdriverout 166.7e-3
rj1453 n8__i5__i7__i7__net3 n6__i5__i7__i7__net3 1.445
rj1454 n751__i1__i14__net1 n749__i1__i14__net1 125e-3
rj1455 n750__i1__i14__net1 n751__i1__i14__net1 125e-3
rj1456 n598__vss n601__vss 166.7e-3
rj1457 n602__vss n597__vss 166.7e-3
rj1458 n595__vss n603__vss 166.7e-3
rj1459 n604__vss n594__vss 166.7e-3
rj1460 n1037__vddio n1050__vddio 166.7e-3
rj1461 n1051__vddio n1040__vddio 166.7e-3
rj1462 n1041__vddio n1052__vddio 166.7e-3
rj1463 n1053__vddio n1043__vddio 166.7e-3
rj1464 n1044__vddio n1054__vddio 166.7e-3
rj1465 n1055__vddio n1046__vddio 166.7e-3
rj1466 n1047__vddio n1056__vddio 166.7e-3
rj1467 n7__i5__i6__net31 n25__i5__i6__net31 1.4217
rj1468 n25__i5__i6__net31 n17__i5__i6__net31 111.9e-3
rj1469 n25__i5__i6__net31 n22__i5__i6__net31 28.86e-3
rj1470 n35__i5__clk_buf n36__i5__clk_buf 500e-3
rj1471 n755__i1__i14__net1 n753__i1__i14__net1 125e-3
rj1472 n754__i1__i14__net1 n755__i1__i14__net1 125e-3
rj1473 n9__i5__i6__i2__net24 n6__i5__i6__i2__net24 176.5e-3
rj1474 n6__i5__i6__i2__net24 n3__i5__i6__i2__net24 178.9e-3
rj1475 n6__i5__i6__i2__net23 n9__i5__i6__i2__net23 489.6e-3
rj1476 n9__i5__i6__i2__net23 n2__i5__i6__i2__net23 236.9e-3
rj1477 n9__i5__i6__i2__net23 n3__i5__i6__i2__net23 278.9e-3
rj1478 n1812__chipdriverout n1813__chipdriverout 166.7e-3
rj1479 n1814__chipdriverout n1815__chipdriverout 166.7e-3
rj1480 n1816__chipdriverout n1817__chipdriverout 166.7e-3
rj1481 n1818__chipdriverout n1819__chipdriverout 166.7e-3
rj1482 n1820__chipdriverout n1821__chipdriverout 166.7e-3
rj1483 n1829__chipdriverout n1843__chipdriverout 166.7e-3
rj1484 n1844__chipdriverout n1832__chipdriverout 166.7e-3
rj1485 n1833__chipdriverout n1845__chipdriverout 166.7e-3
rj1486 n1846__chipdriverout n1835__chipdriverout 166.7e-3
rj1487 n1836__chipdriverout n1847__chipdriverout 166.7e-3
rj1488 n1848__chipdriverout n1838__chipdriverout 166.7e-3
rj1489 n1839__chipdriverout n1849__chipdriverout 166.7e-3
rj1490 n1850__chipdriverout n1841__chipdriverout 166.7e-3
rj1491 n8__i5__r2 n9__i5__r2 250e-3
rj1492 n757__i1__i14__net1 n686__i1__i14__net1 250e-3
rj1493 n688__i1__i14__net1 n757__i1__i14__net1 250e-3
rj1494 n41__reset n40__reset 250e-3
rj1495 n611__vss n614__vss 166.7e-3
rj1496 n615__vss n610__vss 166.7e-3
rj1497 n608__vss n616__vss 166.7e-3
rj1498 n617__vss n607__vss 166.7e-3
rj1499 n1058__vddio n1071__vddio 166.7e-3
rj1500 n1072__vddio n1061__vddio 166.7e-3
rj1501 n1062__vddio n1073__vddio 166.7e-3
rj1502 n1074__vddio n1064__vddio 166.7e-3
rj1503 n1065__vddio n1075__vddio 166.7e-3
rj1504 n1076__vddio n1067__vddio 166.7e-3
rj1505 n1068__vddio n1077__vddio 166.7e-3
rj1506 n690__i1__i14__net1 n762__i1__i14__net1 250e-3
rj1507 n762__i1__i14__net1 n692__i1__i14__net1 250e-3
rj1508 n9__clk_out n8__clk_out 250e-3
rj1509 n1869__chipdriverout n1877__chipdriverout 166.7e-3
rj1510 n1878__chipdriverout n1870__chipdriverout 166.7e-3
rj1511 n1872__chipdriverout n1879__chipdriverout 166.7e-3
rj1512 n1880__chipdriverout n1873__chipdriverout 166.7e-3
rj1513 n1875__chipdriverout n1881__chipdriverout 166.7e-3
rj1514 n1882__chipdriverout n1852__chipdriverout 166.7e-3
rj1515 n1855__chipdriverout n1883__chipdriverout 166.7e-3
rj1516 n1884__chipdriverout n1856__chipdriverout 166.7e-3
rj1517 n1858__chipdriverout n1885__chipdriverout 166.7e-3
rj1518 n1886__chipdriverout n1859__chipdriverout 166.7e-3
rj1519 n1861__chipdriverout n1887__chipdriverout 166.7e-3
rj1520 n1888__chipdriverout n1862__chipdriverout 166.7e-3
rj1521 n1864__chipdriverout n1889__chipdriverout 166.7e-3
rj1522 n765__i1__i14__net1 n767__i1__i14__net1 125e-3
rj1523 n767__i1__i14__net1 n766__i1__i14__net1 125e-3
rj1524 n627__vss n624__vss 166.7e-3
rj1525 n623__vss n628__vss 166.7e-3
rj1526 n629__vss n621__vss 166.7e-3
rj1527 n620__vss n630__vss 166.7e-3
rj1528 n1092__vddio n1079__vddio 166.7e-3
rj1529 n1082__vddio n1093__vddio 166.7e-3
rj1530 n1094__vddio n1083__vddio 166.7e-3
rj1531 n1085__vddio n1095__vddio 166.7e-3
rj1532 n1096__vddio n1086__vddio 166.7e-3
rj1533 n1088__vddio n1097__vddio 166.7e-3
rj1534 n1098__vddio n1089__vddio 166.7e-3
rj1535 n769__i1__i14__net1 n771__i1__i14__net1 125e-3
rj1536 n771__i1__i14__net1 n770__i1__i14__net1 125e-3
rj1537 n632__vss n633__vss 460.8e-3
rj1538 n151__vdd n154__vdd 818.8e-3
rj1539 n1908__chipdriverout n1916__chipdriverout 166.7e-3
rj1540 n1917__chipdriverout n1909__chipdriverout 166.7e-3
rj1541 n1911__chipdriverout n1918__chipdriverout 166.7e-3
rj1542 n1919__chipdriverout n1912__chipdriverout 166.7e-3
rj1543 n1914__chipdriverout n1920__chipdriverout 166.7e-3
rj1544 n1921__chipdriverout n1891__chipdriverout 166.7e-3
rj1545 n1894__chipdriverout n1922__chipdriverout 166.7e-3
rj1546 n1923__chipdriverout n1895__chipdriverout 166.7e-3
rj1547 n1897__chipdriverout n1924__chipdriverout 166.7e-3
rj1548 n1925__chipdriverout n1898__chipdriverout 166.7e-3
rj1549 n1900__chipdriverout n1926__chipdriverout 166.7e-3
rj1550 n1927__chipdriverout n1901__chipdriverout 166.7e-3
rj1551 n1903__chipdriverout n1928__chipdriverout 166.7e-3
rj1552 n775__i1__i14__net1 n773__i1__i14__net1 125e-3
rj1553 n774__i1__i14__net1 n775__i1__i14__net1 125e-3
rj1554 n634__vss n645__vss 509.2e-3
rj1555 n646__vss n642__vss 166.7e-3
rj1556 n641__vss n647__vss 166.7e-3
rj1557 n648__vss n639__vss 166.7e-3
rj1558 n638__vss n649__vss 166.7e-3
rj1559 n1113__vddio n1100__vddio 166.7e-3
rj1560 n1103__vddio n1114__vddio 166.7e-3
rj1561 n1115__vddio n1104__vddio 166.7e-3
rj1562 n1106__vddio n1116__vddio 166.7e-3
rj1563 n1117__vddio n1107__vddio 166.7e-3
rj1564 n1109__vddio n1118__vddio 166.7e-3
rj1565 n1119__vddio n1110__vddio 166.7e-3
rj1566 n157__vdd n158__vdd 566.4e-3
rj1567 n8__i5__i6__net32 n2__i5__i6__net32 1.3485
rj1568 n28__shift n29__shift 1.0669
rj1569 n29__shift n26__shift 28.1e-3
rj1570 n22__shift n29__shift 500e-3
rj1571 n159__vdd n160__vdd 843.7e-3
rj1572 n701__vss n702__vss 723.1e-3
rj1573 n11__i5__r1 n16__i5__r1 166.7e-3
rj1574 n43__i5__clk_buf n44__i5__clk_buf 500e-3
rj1575 n15__i5__i6__net33 n9__i5__i6__net33 838.1e-3
rj1576 n51__i5__clk_buf n52__i5__clk_buf 500e-3
rj1577 n9__i5__i6__i4__net25 n6__i5__i6__i4__net25 176.5e-3
rj1578 n6__i5__i6__i4__net25 n3__i5__i6__i4__net25 178.9e-3
rj1579 n6__i5__i6__i4__net21 n9__i5__i6__i4__net21 494e-3
rj1580 n9__i5__i6__i4__net21 n2__i5__i6__i4__net21 236.9e-3
rj1581 n9__i5__i6__i4__net21 n3__i5__i6__i4__net21 278.9e-3
rj1582 n8__i5__i8__net1 n9__i5__i8__net1 500e-3
rj1583 n712__vss n709__vss 166.7e-3
rj1584 n708__vss n713__vss 166.7e-3
rj1585 n714__vss n706__vss 166.7e-3
rj1586 n705__vss n715__vss 166.7e-3
rj1587 n1187__vddio n1174__vddio 166.7e-3
rj1588 n1177__vddio n1188__vddio 166.7e-3
rj1589 n1189__vddio n1178__vddio 166.7e-3
rj1590 n1180__vddio n1190__vddio 166.7e-3
rj1591 n1191__vddio n1181__vddio 166.7e-3
rj1592 n1183__vddio n1192__vddio 166.7e-3
rj1593 n1193__vddio n1184__vddio 166.7e-3
rj1594 n61__i1__net2 n63__i1__net2 125e-3
rj1595 n63__i1__net2 n62__i1__net2 125e-3
rj1596 n56__i5__clk_buf n57__i5__clk_buf 500e-3
rj1597 n794__i1__i14__net1 n817__i1__i14__net1 166.7e-3
rj1598 n818__i1__i14__net1 n795__i1__i14__net1 166.7e-3
rj1599 n797__i1__i14__net1 n819__i1__i14__net1 166.7e-3
rj1600 n820__i1__i14__net1 n798__i1__i14__net1 166.7e-3
rj1601 n800__i1__i14__net1 n821__i1__i14__net1 166.7e-3
rj1602 n822__i1__i14__net1 n803__i1__i14__net1 166.7e-3
rj1603 n806__i1__i14__net1 n823__i1__i14__net1 166.7e-3
rj1604 n824__i1__i14__net1 n807__i1__i14__net1 166.7e-3
rj1605 n809__i1__i14__net1 n825__i1__i14__net1 166.7e-3
rj1606 n826__i1__i14__net1 n810__i1__i14__net1 166.7e-3
rj1607 n812__i1__i14__net1 n827__i1__i14__net1 166.7e-3
rj1608 n828__i1__i14__net1 n813__i1__i14__net1 166.7e-3
rj1609 n815__i1__i14__net1 n829__i1__i14__net1 166.7e-3
rj1610 n9__i5__i8__i9__net25 n6__i5__i8__i9__net25 176.5e-3
rj1611 n6__i5__i8__i9__net25 n3__i5__i8__i9__net25 178.9e-3
rj1612 n6__i5__i8__i9__net21 n9__i5__i8__i9__net21 494e-3
rj1613 n9__i5__i8__i9__net21 n2__i5__i8__i9__net21 236.9e-3
rj1614 n9__i5__i8__i9__net21 n3__i5__i8__i9__net21 278.9e-3
rj1615 n69__i1__net2 n71__i1__net2 125e-3
rj1616 n71__i1__net2 n70__i1__net2 125e-3
rj1617 n28__i5__i6__net31 n37__i5__i6__net31 1.4217
rj1618 n37__i5__i6__net31 n29__i5__i6__net31 111.9e-3
rj1619 n37__i5__i6__net31 n30__i5__i6__net31 28.86e-3
rj1620 n725__vss n722__vss 166.7e-3
rj1621 n721__vss n726__vss 166.7e-3
rj1622 n727__vss n719__vss 166.7e-3
rj1623 n718__vss n728__vss 166.7e-3
rj1624 n1214__vddio n1201__vddio 166.7e-3
rj1625 n1204__vddio n1215__vddio 166.7e-3
rj1626 n1216__vddio n1205__vddio 166.7e-3
rj1627 n1207__vddio n1217__vddio 166.7e-3
rj1628 n1218__vddio n1208__vddio 166.7e-3
rj1629 n1210__vddio n1219__vddio 166.7e-3
rj1630 n1220__vddio n1211__vddio 166.7e-3
rj1631 n58__i5__clk_buf n59__i5__clk_buf 500e-3
rj1632 n79__i1__net2 n77__i1__net2 125e-3
rj1633 n78__i1__net2 n79__i1__net2 125e-3
rj1634 n9__i5__i6__i4__net24 n6__i5__i6__i4__net24 176.5e-3
rj1635 n6__i5__i6__i4__net24 n3__i5__i6__i4__net24 178.9e-3
rj1636 n6__i5__i6__i4__net23 n9__i5__i6__i4__net23 489.6e-3
rj1637 n9__i5__i6__i4__net23 n2__i5__i6__i4__net23 236.9e-3
rj1638 n9__i5__i6__i4__net23 n3__i5__i6__i4__net23 278.9e-3
rj1639 n833__i1__i14__net1 n856__i1__i14__net1 166.7e-3
rj1640 n857__i1__i14__net1 n834__i1__i14__net1 166.7e-3
rj1641 n836__i1__i14__net1 n858__i1__i14__net1 166.7e-3
rj1642 n859__i1__i14__net1 n837__i1__i14__net1 166.7e-3
rj1643 n839__i1__i14__net1 n860__i1__i14__net1 166.7e-3
rj1644 n861__i1__i14__net1 n842__i1__i14__net1 166.7e-3
rj1645 n845__i1__i14__net1 n862__i1__i14__net1 166.7e-3
rj1646 n863__i1__i14__net1 n846__i1__i14__net1 166.7e-3
rj1647 n848__i1__i14__net1 n864__i1__i14__net1 166.7e-3
rj1648 n865__i1__i14__net1 n849__i1__i14__net1 166.7e-3
rj1649 n851__i1__i14__net1 n866__i1__i14__net1 166.7e-3
rj1650 n867__i1__i14__net1 n852__i1__i14__net1 166.7e-3
rj1651 n854__i1__i14__net1 n868__i1__i14__net1 166.7e-3
rj1652 n45__reset n51__reset 250e-3
rj1653 n14__i1__net2 n82__i1__net2 250e-3
rj1654 n82__i1__net2 n16__i1__net2 250e-3
rj1655 n7__i5__i8__net4 n17__i5__i8__net4 1.1119
rj1656 n17__i5__i8__net4 n12__i5__i8__net4 1.0819
rj1657 n17__i5__i8__net4 n15__i5__i8__net4 422.2e-3
rj1658 n735__vss n738__vss 166.7e-3
rj1659 n739__vss n734__vss 166.7e-3
rj1660 n732__vss n740__vss 166.7e-3
rj1661 n741__vss n731__vss 166.7e-3
rj1662 n1222__vddio n1235__vddio 166.7e-3
rj1663 n1236__vddio n1225__vddio 166.7e-3
rj1664 n1226__vddio n1237__vddio 166.7e-3
rj1665 n1238__vddio n1228__vddio 166.7e-3
rj1666 n1229__vddio n1239__vddio 166.7e-3
rj1667 n1240__vddio n1231__vddio 166.7e-3
rj1668 n1232__vddio n1241__vddio 166.7e-3
rj1669 n63__i5__clk_buf n64__i5__clk_buf 500e-3
rj1670 n91__i1__net2 n89__i1__net2 125e-3
rj1671 n90__i1__net2 n91__i1__net2 125e-3
rj1672 n7__i5__i8__i9__net24 n6__i5__i8__i9__net24 426.5e-3
rj1673 n6__i5__i8__i9__net24 n3__i5__i8__i9__net24 178.9e-3
rj1674 n6__i5__i8__i9__net23 n7__i5__i8__i9__net23 489.6e-3
rj1675 n7__i5__i8__i9__net23 n2__i5__i8__i9__net23 236.9e-3
rj1676 n7__i5__i8__i9__net23 n3__i5__i8__i9__net23 278.9e-3
rj1677 n895__i1__i14__net1 n872__i1__i14__net1 166.7e-3
rj1678 n873__i1__i14__net1 n896__i1__i14__net1 166.7e-3
rj1679 n897__i1__i14__net1 n875__i1__i14__net1 166.7e-3
rj1680 n876__i1__i14__net1 n898__i1__i14__net1 166.7e-3
rj1681 n899__i1__i14__net1 n878__i1__i14__net1 166.7e-3
rj1682 n881__i1__i14__net1 n900__i1__i14__net1 166.7e-3
rj1683 n901__i1__i14__net1 n884__i1__i14__net1 166.7e-3
rj1684 n885__i1__i14__net1 n902__i1__i14__net1 166.7e-3
rj1685 n903__i1__i14__net1 n887__i1__i14__net1 166.7e-3
rj1686 n888__i1__i14__net1 n904__i1__i14__net1 166.7e-3
rj1687 n905__i1__i14__net1 n890__i1__i14__net1 166.7e-3
rj1688 n891__i1__i14__net1 n906__i1__i14__net1 166.7e-3
rj1689 n907__i1__i14__net1 n893__i1__i14__net1 166.7e-3
rj1690 n99__i1__net2 n97__i1__net2 125e-3
rj1691 n98__i1__net2 n99__i1__net2 125e-3
rj1692 n54__reset n55__reset 250e-3
rj1693 n742__vss n743__vss 166.7e-3
rj1694 n744__vss n745__vss 166.7e-3
rj1695 n746__vss n747__vss 166.7e-3
rj1696 n748__vss n749__vss 166.7e-3
rj1697 n1242__vddio n1243__vddio 166.7e-3
rj1698 n1244__vddio n1245__vddio 166.7e-3
rj1699 n1246__vddio n1247__vddio 166.7e-3
rj1700 n1248__vddio n1249__vddio 166.7e-3
rj1701 n1250__vddio n1251__vddio 166.7e-3
rj1702 n1252__vddio n1253__vddio 166.7e-3
rj1703 n1254__vddio n1255__vddio 166.7e-3
rj1704 n109__i1__net2 n111__i1__net2 125e-3
rj1705 n111__i1__net2 n110__i1__net2 125e-3
rj1706 n911__i1__i14__net1 n934__i1__i14__net1 166.7e-3
rj1707 n935__i1__i14__net1 n912__i1__i14__net1 166.7e-3
rj1708 n914__i1__i14__net1 n936__i1__i14__net1 166.7e-3
rj1709 n937__i1__i14__net1 n915__i1__i14__net1 166.7e-3
rj1710 n917__i1__i14__net1 n938__i1__i14__net1 166.7e-3
rj1711 n939__i1__i14__net1 n920__i1__i14__net1 166.7e-3
rj1712 n923__i1__i14__net1 n940__i1__i14__net1 166.7e-3
rj1713 n941__i1__i14__net1 n924__i1__i14__net1 166.7e-3
rj1714 n926__i1__i14__net1 n942__i1__i14__net1 166.7e-3
rj1715 n943__i1__i14__net1 n927__i1__i14__net1 166.7e-3
rj1716 n929__i1__i14__net1 n944__i1__i14__net1 166.7e-3
rj1717 n945__i1__i14__net1 n930__i1__i14__net1 166.7e-3
rj1718 n932__i1__i14__net1 n946__i1__i14__net1 166.7e-3
rj1719 n117__i1__net2 n30__i1__net2 250e-3
rj1720 n32__i1__net2 n117__i1__net2 250e-3
rj1721 n8__i5__i6__net34 n2__i5__i6__net34 1.3504
rj1722 n16__i5__i8__net2 n17__i5__i8__net2 500e-3
rj1723 n764__vss n761__vss 166.7e-3
rj1724 n760__vss n765__vss 166.7e-3
rj1725 n766__vss n758__vss 166.7e-3
rj1726 n757__vss n767__vss 166.7e-3
rj1727 n1277__vddio n1264__vddio 166.7e-3
rj1728 n1267__vddio n1278__vddio 166.7e-3
rj1729 n1279__vddio n1268__vddio 166.7e-3
rj1730 n1270__vddio n1280__vddio 166.7e-3
rj1731 n1281__vddio n1271__vddio 166.7e-3
rj1732 n1273__vddio n1282__vddio 166.7e-3
rj1733 n1283__vddio n1274__vddio 166.7e-3
rj1734 n38__shift n39__shift 1.0669
rj1735 n39__shift n36__shift 28.1e-3
rj1736 n35__shift n39__shift 500e-3
rj1737 n125__i1__net2 n34__i1__net2 250e-3
rj1738 n36__i1__net2 n125__i1__net2 250e-3
rj1739 n950__i1__i14__net1 n973__i1__i14__net1 166.7e-3
rj1740 n974__i1__i14__net1 n951__i1__i14__net1 166.7e-3
rj1741 n953__i1__i14__net1 n975__i1__i14__net1 166.7e-3
rj1742 n976__i1__i14__net1 n954__i1__i14__net1 166.7e-3
rj1743 n956__i1__i14__net1 n977__i1__i14__net1 166.7e-3
rj1744 n978__i1__i14__net1 n959__i1__i14__net1 166.7e-3
rj1745 n962__i1__i14__net1 n979__i1__i14__net1 166.7e-3
rj1746 n980__i1__i14__net1 n963__i1__i14__net1 166.7e-3
rj1747 n965__i1__i14__net1 n981__i1__i14__net1 166.7e-3
rj1748 n982__i1__i14__net1 n966__i1__i14__net1 166.7e-3
rj1749 n968__i1__i14__net1 n983__i1__i14__net1 166.7e-3
rj1750 n984__i1__i14__net1 n969__i1__i14__net1 166.7e-3
rj1751 n971__i1__i14__net1 n985__i1__i14__net1 166.7e-3
rj1752 n129__i1__net2 n131__i1__net2 125e-3
rj1753 n131__i1__net2 n130__i1__net2 125e-3
rj1754 n12__i5__r0 n14__i5__r0 333.3e-3
rj1755 n774__vss n777__vss 166.7e-3
rj1756 n778__vss n773__vss 166.7e-3
rj1757 n771__vss n779__vss 166.7e-3
rj1758 n780__vss n770__vss 166.7e-3
rj1759 n1295__vddio n1308__vddio 166.7e-3
rj1760 n1309__vddio n1298__vddio 166.7e-3
rj1761 n1299__vddio n1310__vddio 166.7e-3
rj1762 n1311__vddio n1301__vddio 166.7e-3
rj1763 n1302__vddio n1312__vddio 166.7e-3
rj1764 n1313__vddio n1304__vddio 166.7e-3
rj1765 n1305__vddio n1314__vddio 166.7e-3
rj1766 n141__i1__net2 n143__i1__net2 125e-3
rj1767 n143__i1__net2 n142__i1__net2 125e-3
rj1768 n989__i1__i14__net1 n1012__i1__i14__net1 166.7e-3
rj1769 n1013__i1__i14__net1 n990__i1__i14__net1 166.7e-3
rj1770 n992__i1__i14__net1 n1014__i1__i14__net1 166.7e-3
rj1771 n1015__i1__i14__net1 n993__i1__i14__net1 166.7e-3
rj1772 n995__i1__i14__net1 n1016__i1__i14__net1 166.7e-3
rj1773 n1017__i1__i14__net1 n998__i1__i14__net1 166.7e-3
rj1774 n1001__i1__i14__net1 n1018__i1__i14__net1 166.7e-3
rj1775 n1019__i1__i14__net1 n1002__i1__i14__net1 166.7e-3
rj1776 n1004__i1__i14__net1 n1020__i1__i14__net1 166.7e-3
rj1777 n1021__i1__i14__net1 n1005__i1__i14__net1 166.7e-3
rj1778 n1007__i1__i14__net1 n1022__i1__i14__net1 166.7e-3
rj1779 n1023__i1__i14__net1 n1008__i1__i14__net1 166.7e-3
rj1780 n1010__i1__i14__net1 n1024__i1__i14__net1 166.7e-3
rj1781 n15__i5__i6__net35 n9__i5__i6__net35 838.1e-3
rj1782 n151__i1__net2 n149__i1__net2 125e-3
rj1783 n150__i1__net2 n151__i1__net2 125e-3
rj1784 n790__vss n787__vss 166.7e-3
rj1785 n786__vss n791__vss 166.7e-3
rj1786 n792__vss n784__vss 166.7e-3
rj1787 n783__vss n793__vss 166.7e-3
rj1788 n1329__vddio n1316__vddio 166.7e-3
rj1789 n1319__vddio n1330__vddio 166.7e-3
rj1790 n1331__vddio n1320__vddio 166.7e-3
rj1791 n1322__vddio n1332__vddio 166.7e-3
rj1792 n1333__vddio n1323__vddio 166.7e-3
rj1793 n1325__vddio n1334__vddio 166.7e-3
rj1794 n1335__vddio n1326__vddio 166.7e-3
rj1795 n9__i5__i8__net5 n8__i5__i8__net5 250e-3
rj1796 n159__i1__net2 n157__i1__net2 125e-3
rj1797 n158__i1__net2 n159__i1__net2 125e-3
rj1798 n65__i5__clk_buf n66__i5__clk_buf 500e-3
rj1799 n1043__i1__i14__net1 n1051__i1__i14__net1 166.7e-3
rj1800 n1052__i1__i14__net1 n1044__i1__i14__net1 166.7e-3
rj1801 n1046__i1__i14__net1 n1053__i1__i14__net1 166.7e-3
rj1802 n1054__i1__i14__net1 n1047__i1__i14__net1 166.7e-3
rj1803 n1049__i1__i14__net1 n1055__i1__i14__net1 166.7e-3
rj1804 n1056__i1__i14__net1 n1026__i1__i14__net1 166.7e-3
rj1805 n1029__i1__i14__net1 n1057__i1__i14__net1 166.7e-3
rj1806 n1058__i1__i14__net1 n1030__i1__i14__net1 166.7e-3
rj1807 n1032__i1__i14__net1 n1059__i1__i14__net1 166.7e-3
rj1808 n1060__i1__i14__net1 n1033__i1__i14__net1 166.7e-3
rj1809 n1035__i1__i14__net1 n1061__i1__i14__net1 166.7e-3
rj1810 n1062__i1__i14__net1 n1036__i1__i14__net1 166.7e-3
rj1811 n1038__i1__i14__net1 n1063__i1__i14__net1 166.7e-3
rj1813 n33__i5__i8__net2 n27__i5__i8__net2 1.0556
rj1814 n161__i1__net2 n54__i1__net2 250e-3
rj1815 n56__i1__net2 n161__i1__net2 250e-3
rj1816 n7__i5__i6__i5__net25 n6__i5__i6__i5__net25 426.5e-3
rj1817 n6__i5__i6__i5__net25 n3__i5__i6__i5__net25 178.9e-3
rj1818 n6__i5__i6__i5__net21 n7__i5__i6__i5__net21 494e-3
rj1819 n7__i5__i6__i5__net21 n2__i5__i6__i5__net21 236.9e-3
rj1820 n7__i5__i6__i5__net21 n3__i5__i6__i5__net21 278.9e-3
rj1821 n7__i5__i8__i10__net25 n6__i5__i8__i10__net25 426.5e-3
rj1822 n6__i5__i8__i10__net25 n3__i5__i8__i10__net25 178.9e-3
rj1823 n6__i5__i8__i10__net21 n7__i5__i8__i10__net21 494e-3
rj1824 n7__i5__i8__i10__net21 n2__i5__i8__i10__net21 254.9e-3
rj1825 n7__i5__i8__i10__net21 n3__i5__i8__i10__net21 278.9e-3
rj1826 n794__vss n795__vss 166.7e-3
rj1827 n796__vss n797__vss 166.7e-3
rj1828 n798__vss n799__vss 166.7e-3
rj1829 n800__vss n801__vss 166.7e-3
rj1830 n1336__vddio n1337__vddio 166.7e-3
rj1831 n1338__vddio n1339__vddio 166.7e-3
rj1832 n1340__vddio n1341__vddio 166.7e-3
rj1833 n1342__vddio n1343__vddio 166.7e-3
rj1834 n1344__vddio n1345__vddio 166.7e-3
rj1835 n1346__vddio n1347__vddio 166.7e-3
rj1836 n1348__vddio n1349__vddio 166.7e-3
rj1837 n165__i1__net2 n58__i1__net2 250e-3
rj1838 n60__i1__net2 n165__i1__net2 250e-3
rj1839 n1064__i1__i14__net1 n1065__i1__i14__net1 166.7e-3
rj1840 n1066__i1__i14__net1 n1067__i1__i14__net1 166.7e-3
rj1841 n1068__i1__i14__net1 n1069__i1__i14__net1 166.7e-3
rj1842 n1070__i1__i14__net1 n1071__i1__i14__net1 166.7e-3
rj1843 n1072__i1__i14__net1 n1073__i1__i14__net1 166.7e-3
rj1844 n1074__i1__i14__net1 n1075__i1__i14__net1 166.7e-3
rj1845 n1076__i1__i14__net1 n1077__i1__i14__net1 166.7e-3
rj1846 n1078__i1__i14__net1 n1079__i1__i14__net1 166.7e-3
rj1847 n1080__i1__i14__net1 n1081__i1__i14__net1 166.7e-3
rj1848 n1082__i1__i14__net1 n1083__i1__i14__net1 166.7e-3
rj1849 n1084__i1__i14__net1 n1085__i1__i14__net1 166.7e-3
rj1850 n1086__i1__i14__net1 n1087__i1__i14__net1 166.7e-3
rj1851 n1088__i1__i14__net1 n1089__i1__i14__net1 166.7e-3
rj1852 n173__i1__net2 n169__i1__net2 125e-3
rj1853 n170__i1__net2 n173__i1__net2 125e-3
rj1854 n816__vss n813__vss 166.7e-3
rj1855 n812__vss n817__vss 166.7e-3
rj1856 n818__vss n810__vss 166.7e-3
rj1857 n809__vss n819__vss 166.7e-3
rj1858 n1371__vddio n1358__vddio 166.7e-3
rj1859 n1361__vddio n1372__vddio 166.7e-3
rj1860 n1373__vddio n1362__vddio 166.7e-3
rj1861 n1364__vddio n1374__vddio 166.7e-3
rj1862 n1375__vddio n1365__vddio 166.7e-3
rj1863 n1367__vddio n1376__vddio 166.7e-3
rj1864 n1377__vddio n1368__vddio 166.7e-3
rj1865 n44__i5__i6__net31 n45__i5__i6__net31 921.7e-3
rj1866 n45__i5__i6__net31 n41__i5__i6__net31 111.9e-3
rj1867 n45__i5__i6__net31 n42__i5__i6__net31 28.86e-3
rj1868 n27__i5__i8__net1 n26__i5__i8__net1 1.0273
rj1869 n26__i5__i8__net1 n24__i5__i8__net1 467.5e-3
rj1871 n19__i5__i8__net1 n24__i5__i8__net1 250e-3
rj1872 n67__i5__clk_buf n68__i5__clk_buf 500e-3
rj1873 n35__i5__i8__net2 n36__i5__i8__net2 500e-3
rj1874 n175__i1__net2 n171__i1__net2 125e-3
rj1875 n172__i1__net2 n175__i1__net2 125e-3
rj1876 n1106__i1__i14__net1 n1129__i1__i14__net1 166.7e-3
rj1877 n1130__i1__i14__net1 n1107__i1__i14__net1 166.7e-3
rj1878 n1109__i1__i14__net1 n1131__i1__i14__net1 166.7e-3
rj1879 n1132__i1__i14__net1 n1110__i1__i14__net1 166.7e-3
rj1880 n1112__i1__i14__net1 n1133__i1__i14__net1 166.7e-3
rj1881 n1134__i1__i14__net1 n1115__i1__i14__net1 166.7e-3
rj1882 n1118__i1__i14__net1 n1135__i1__i14__net1 166.7e-3
rj1883 n1136__i1__i14__net1 n1119__i1__i14__net1 166.7e-3
rj1884 n1121__i1__i14__net1 n1137__i1__i14__net1 166.7e-3
rj1885 n1138__i1__i14__net1 n1122__i1__i14__net1 166.7e-3
rj1886 n1124__i1__i14__net1 n1139__i1__i14__net1 166.7e-3
rj1887 n1140__i1__i14__net1 n1125__i1__i14__net1 166.7e-3
rj1888 n1127__i1__i14__net1 n1141__i1__i14__net1 166.7e-3
rj1889 n7__i5__i6__i5__net24 n6__i5__i6__i5__net24 426.5e-3
rj1890 n6__i5__i6__i5__net24 n3__i5__i6__i5__net24 178.9e-3
rj1891 n6__i5__i6__i5__net23 n7__i5__i6__i5__net23 489.6e-3
rj1892 n7__i5__i6__i5__net23 n2__i5__i6__i5__net23 236.9e-3
rj1893 n7__i5__i6__i5__net23 n3__i5__i6__i5__net23 278.9e-3
rj1894 n9__i5__i8__i10__net24 n6__i5__i8__i10__net24 176.5e-3
rj1895 n6__i5__i8__i10__net24 n3__i5__i8__i10__net24 178.9e-3
rj1896 n6__i5__i8__i10__net23 n9__i5__i8__i10__net23 489.6e-3
rj1897 n9__i5__i8__i10__net23 n2__i5__i8__i10__net23 236.9e-3
rj1898 n9__i5__i8__i10__net23 n3__i5__i8__i10__net23 278.9e-3
rj1899 n177__i1__net2 n179__i1__net2 125e-3
rj1900 n179__i1__net2 n178__i1__net2 125e-3
rj1901 n68__reset n70__reset 250e-3
rj1902 n69__reset n71__reset 250e-3
rj1903 n826__vss n829__vss 166.7e-3
rj1904 n830__vss n825__vss 166.7e-3
rj1905 n823__vss n831__vss 166.7e-3
rj1906 n832__vss n822__vss 166.7e-3
rj1907 n1379__vddio n1392__vddio 166.7e-3
rj1908 n1393__vddio n1382__vddio 166.7e-3
rj1909 n1383__vddio n1394__vddio 166.7e-3
rj1910 n1395__vddio n1385__vddio 166.7e-3
rj1911 n1386__vddio n1396__vddio 166.7e-3
rj1912 n1397__vddio n1388__vddio 166.7e-3
rj1913 n1389__vddio n1398__vddio 166.7e-3
rj1914 n94__i1__net2 n186__i1__net2 250e-3
rj1915 n186__i1__net2 n96__i1__net2 250e-3
rj1916 n1168__i1__i14__net1 n1145__i1__i14__net1 166.7e-3
rj1917 n1146__i1__i14__net1 n1169__i1__i14__net1 166.7e-3
rj1918 n1170__i1__i14__net1 n1148__i1__i14__net1 166.7e-3
rj1919 n1149__i1__i14__net1 n1171__i1__i14__net1 166.7e-3
rj1920 n1172__i1__i14__net1 n1151__i1__i14__net1 166.7e-3
rj1921 n1154__i1__i14__net1 n1173__i1__i14__net1 166.7e-3
rj1922 n1174__i1__i14__net1 n1157__i1__i14__net1 166.7e-3
rj1923 n1158__i1__i14__net1 n1175__i1__i14__net1 166.7e-3
rj1924 n1176__i1__i14__net1 n1160__i1__i14__net1 166.7e-3
rj1925 n1161__i1__i14__net1 n1177__i1__i14__net1 166.7e-3
rj1926 n1178__i1__i14__net1 n1163__i1__i14__net1 166.7e-3
rj1927 n1164__i1__i14__net1 n1179__i1__i14__net1 166.7e-3
rj1928 n1180__i1__i14__net1 n1166__i1__i14__net1 166.7e-3
rj1929 n191__i1__net2 n189__i1__net2 125e-3
rj1930 n190__i1__net2 n191__i1__net2 125e-3
rj1931 n839__vss n842__vss 166.7e-3
rj1932 n843__vss n838__vss 166.7e-3
rj1933 n836__vss n844__vss 166.7e-3
rj1934 n845__vss n835__vss 166.7e-3
rj1935 n1410__vddio n1423__vddio 166.7e-3
rj1936 n1424__vddio n1413__vddio 166.7e-3
rj1937 n1414__vddio n1425__vddio 166.7e-3
rj1938 n1426__vddio n1416__vddio 166.7e-3
rj1939 n1417__vddio n1427__vddio 166.7e-3
rj1940 n1428__vddio n1419__vddio 166.7e-3
rj1941 n1420__vddio n1429__vddio 166.7e-3
rj1942 n195__i1__net2 n193__i1__net2 125e-3
rj1943 n194__i1__net2 n195__i1__net2 125e-3
rj1944 n1199__i1__i14__net1 n1207__i1__i14__net1 166.7e-3
rj1945 n1208__i1__i14__net1 n1200__i1__i14__net1 166.7e-3
rj1946 n1202__i1__i14__net1 n1209__i1__i14__net1 166.7e-3
rj1947 n1210__i1__i14__net1 n1203__i1__i14__net1 166.7e-3
rj1948 n1205__i1__i14__net1 n1211__i1__i14__net1 166.7e-3
rj1949 n1212__i1__i14__net1 n1182__i1__i14__net1 166.7e-3
rj1950 n1185__i1__i14__net1 n1213__i1__i14__net1 166.7e-3
rj1951 n1214__i1__i14__net1 n1186__i1__i14__net1 166.7e-3
rj1952 n1188__i1__i14__net1 n1215__i1__i14__net1 166.7e-3
rj1953 n1216__i1__i14__net1 n1189__i1__i14__net1 166.7e-3
rj1954 n1191__i1__i14__net1 n1217__i1__i14__net1 166.7e-3
rj1955 n1218__i1__i14__net1 n1192__i1__i14__net1 166.7e-3
rj1956 n1194__i1__i14__net1 n1219__i1__i14__net1 166.7e-3
rj1957 n199__i1__net2 n197__i1__net2 125e-3
rj1958 n198__i1__net2 n199__i1__net2 125e-3
rj1959 n855__vss n852__vss 166.7e-3
rj1960 n851__vss n856__vss 166.7e-3
rj1961 n857__vss n849__vss 166.7e-3
rj1962 n848__vss n858__vss 166.7e-3
rj1963 n1444__vddio n1431__vddio 166.7e-3
rj1964 n1434__vddio n1445__vddio 166.7e-3
rj1965 n1446__vddio n1435__vddio 166.7e-3
rj1966 n1437__vddio n1447__vddio 166.7e-3
rj1967 n1448__vddio n1438__vddio 166.7e-3
rj1968 n1440__vddio n1449__vddio 166.7e-3
rj1969 n1450__vddio n1441__vddio 166.7e-3
rj1970 n201__i1__net2 n203__i1__net2 125e-3
rj1971 n203__i1__net2 n202__i1__net2 125e-3
rj1972 n11__i5__i8__net5 n12__i5__i8__net5 500e-3
rj1973 n1246__i1__i14__net1 n1238__i1__i14__net1 166.7e-3
rj1974 n1239__i1__i14__net1 n1247__i1__i14__net1 166.7e-3
rj1975 n1248__i1__i14__net1 n1241__i1__i14__net1 166.7e-3
rj1976 n1242__i1__i14__net1 n1249__i1__i14__net1 166.7e-3
rj1977 n1250__i1__i14__net1 n1244__i1__i14__net1 166.7e-3
rj1978 n1221__i1__i14__net1 n1251__i1__i14__net1 166.7e-3
rj1979 n1252__i1__i14__net1 n1224__i1__i14__net1 166.7e-3
rj1980 n1225__i1__i14__net1 n1253__i1__i14__net1 166.7e-3
rj1981 n1254__i1__i14__net1 n1227__i1__i14__net1 166.7e-3
rj1982 n1228__i1__i14__net1 n1255__i1__i14__net1 166.7e-3
rj1983 n1256__i1__i14__net1 n1230__i1__i14__net1 166.7e-3
rj1984 n1231__i1__i14__net1 n1257__i1__i14__net1 166.7e-3
rj1985 n1258__i1__i14__net1 n1233__i1__i14__net1 166.7e-3
rj1986 n205__i1__net2 n207__i1__net2 125e-3
rj1987 n207__i1__net2 n206__i1__net2 125e-3
rj1988 n865__vss n868__vss 166.7e-3
rj1989 n869__vss n864__vss 166.7e-3
rj1990 n862__vss n870__vss 166.7e-3
rj1991 n871__vss n861__vss 166.7e-3
rj1992 n1452__vddio n1465__vddio 166.7e-3
rj1993 n1466__vddio n1455__vddio 166.7e-3
rj1994 n1456__vddio n1467__vddio 166.7e-3
rj1995 n1468__vddio n1458__vddio 166.7e-3
rj1996 n1459__vddio n1469__vddio 166.7e-3
rj1997 n1470__vddio n1461__vddio 166.7e-3
rj1998 n1462__vddio n1471__vddio 166.7e-3
rj1999 n94__i5__clk4 n98__i5__clk4 526.9e-3
rj2000 n98__i5__clk4 n101__i5__clk4 93.78e-3
rj2001 n6__piso_out n18__piso_out 250e-3
rj2002 n209__i1__net2 n211__i1__net2 125e-3
rj2003 n211__i1__net2 n210__i1__net2 125e-3
rj2004 n38__i5__i8__net2 n37__i5__i8__net2 22.62e-3
rj2005 n1285__i1__i14__net1 n1262__i1__i14__net1 166.7e-3
rj2006 n1263__i1__i14__net1 n1286__i1__i14__net1 166.7e-3
rj2007 n1287__i1__i14__net1 n1265__i1__i14__net1 166.7e-3
rj2008 n1266__i1__i14__net1 n1288__i1__i14__net1 166.7e-3
rj2009 n1289__i1__i14__net1 n1268__i1__i14__net1 166.7e-3
rj2010 n1271__i1__i14__net1 n1290__i1__i14__net1 166.7e-3
rj2011 n1291__i1__i14__net1 n1274__i1__i14__net1 166.7e-3
rj2012 n1275__i1__i14__net1 n1292__i1__i14__net1 166.7e-3
rj2013 n1293__i1__i14__net1 n1277__i1__i14__net1 166.7e-3
rj2014 n1278__i1__i14__net1 n1294__i1__i14__net1 166.7e-3
rj2015 n1295__i1__i14__net1 n1280__i1__i14__net1 166.7e-3
rj2016 n1281__i1__i14__net1 n1296__i1__i14__net1 166.7e-3
rj2017 n1297__i1__i14__net1 n1283__i1__i14__net1 166.7e-3
rj2018 n213__i1__net2 n146__i1__net2 250e-3
rj2019 n148__i1__net2 n213__i1__net2 250e-3
rj2020 n872__vss n873__vss 166.7e-3
rj2021 n874__vss n875__vss 166.7e-3
rj2022 n876__vss n877__vss 166.7e-3
rj2023 n878__vss n879__vss 166.7e-3
rj2024 n1472__vddio n1473__vddio 166.7e-3
rj2025 n1474__vddio n1475__vddio 166.7e-3
rj2026 n1476__vddio n1477__vddio 166.7e-3
rj2027 n1478__vddio n1479__vddio 166.7e-3
rj2028 n1480__vddio n1481__vddio 166.7e-3
rj2029 n1482__vddio n1483__vddio 166.7e-3
rj2030 n1484__vddio n1485__vddio 166.7e-3
rj2031 piso_outinv n2__piso_outinv 500e-3
rj2032 n219__i1__net2 n217__i1__net2 125e-3
rj2033 n218__i1__net2 n219__i1__net2 125e-3
rj2034 n1298__i1__i14__net1 n1299__i1__i14__net1 166.7e-3
rj2035 n1300__i1__i14__net1 n1301__i1__i14__net1 166.7e-3
rj2036 n1302__i1__i14__net1 n1303__i1__i14__net1 166.7e-3
rj2037 n1304__i1__i14__net1 n1305__i1__i14__net1 166.7e-3
rj2038 n1306__i1__i14__net1 n1307__i1__i14__net1 166.7e-3
rj2039 n1308__i1__i14__net1 n1309__i1__i14__net1 166.7e-3
rj2040 n1310__i1__i14__net1 n1311__i1__i14__net1 166.7e-3
rj2041 n1312__i1__i14__net1 n1313__i1__i14__net1 166.7e-3
rj2042 n1314__i1__i14__net1 n1315__i1__i14__net1 166.7e-3
rj2043 n1316__i1__i14__net1 n1317__i1__i14__net1 166.7e-3
rj2044 n1318__i1__i14__net1 n1319__i1__i14__net1 166.7e-3
rj2045 n1320__i1__i14__net1 n1321__i1__i14__net1 166.7e-3
rj2046 n1322__i1__i14__net1 n1323__i1__i14__net1 166.7e-3
rj2047 n221__i1__net2 n223__i1__net2 125e-3
rj2048 n223__i1__net2 n222__i1__net2 125e-3
rj2049 n40__shift shift 633.2e-3
rj2050 shift n45__shift 638.5e-3
rj2051 n885__vss n886__vss 166.7e-3
rj2052 n887__vss n888__vss 166.7e-3
rj2053 n889__vss n890__vss 166.7e-3
rj2054 n891__vss n892__vss 166.7e-3
rj2055 n1493__vddio n1494__vddio 166.7e-3
rj2056 n1495__vddio n1496__vddio 166.7e-3
rj2057 n1497__vddio n1498__vddio 166.7e-3
rj2058 n1499__vddio n1500__vddio 166.7e-3
rj2059 n1501__vddio n1502__vddio 166.7e-3
rj2060 n1503__vddio n1504__vddio 166.7e-3
rj2061 n1505__vddio n1506__vddio 166.7e-3
rj2063 n376__vdd n378__vdd 440.7e-3
rj2065 n378__vdd n380__vdd 440.7e-3
rj2067 n380__vdd n382__vdd 440.7e-3
rj2069 n382__vdd n384__vdd 440.7e-3
rj2070 n384__vdd n154__vdd 12.5e-3
rj2071 n184__vdd n376__vdd 12.5e-3
rj2072 n189__vdd n378__vdd 12.5e-3
rj2073 n194__vdd n380__vdd 12.5e-3
rj2074 n198__vdd n382__vdd 12.5e-3
rj2076 n893__vss n913__vss 147.4e-3
rj2078 n913__vss n884__vss 114.4e-3
rj2080 n913__vss n916__vss 90.27e-3
rj2081 n916__vss n867__vss 95.53e-3
rj2082 n867__vss n895__vss 83.33e-3
rj2083 n916__vss n917__vss 65.33e-3
rj2084 n917__vss n854__vss 95.53e-3
rj2086 n917__vss n919__vss 49.2e-3
rj2088 n919__vss n841__vss 114.4e-3
rj2089 n841__vss n897__vss 83.33e-3
rj2090 n919__vss n921__vss 86.26e-3
rj2091 n921__vss n828__vss 95.53e-3
rj2093 n921__vss n923__vss 70.34e-3
rj2094 n923__vss n815__vss 95.53e-3
rj2096 n923__vss n925__vss 65.33e-3
rj2097 n925__vss n806__vss 95.53e-3
rj2098 n806__vss n900__vss 83.33e-3
rj2099 n925__vss n926__vss 50.2e-3
rj2101 n926__vss n789__vss 114.4e-3
rj2102 n789__vss n901__vss 83.33e-3
rj2103 n926__vss n928__vss 85.26e-3
rj2104 n928__vss n776__vss 95.53e-3
rj2106 n928__vss n930__vss 70.34e-3
rj2107 n930__vss n763__vss 95.53e-3
rj2109 n930__vss n932__vss 65.33e-3
rj2110 n932__vss n754__vss 95.53e-3
rj2112 n932__vss n934__vss 51.2e-3
rj2114 n934__vss n737__vss 114.4e-3
rj2116 n934__vss n937__vss 84.26e-3
rj2117 n937__vss n724__vss 95.53e-3
rj2118 n724__vss n906__vss 83.33e-3
rj2119 n937__vss n938__vss 70.34e-3
rj2120 n938__vss n711__vss 95.53e-3
rj2122 n938__vss n939__vss 120.3e-3
rj2124 n939__vss n941__vss 105.3e-3
rj2125 n941__vss n644__vss 95.53e-3
rj2127 n941__vss n942__vss 65.33e-3
rj2128 n942__vss n626__vss 95.53e-3
rj2130 n942__vss n944__vss 104.3e-3
rj2132 n944__vss n613__vss 114.4e-3
rj2134 n944__vss n600__vss 114.4e-3
rj2135 n600__vss n653__vss 83.33e-3
rj2136 n944__vss n947__vss 104.3e-3
rj2137 n947__vss n591__vss 95.53e-3
rj2138 n591__vss n654__vss 83.33e-3
rj2139 n947__vss n948__vss 65.33e-3
rj2140 n948__vss n574__vss 95.53e-3
rj2141 n574__vss n655__vss 83.33e-3
rj2142 n948__vss n949__vss 105.3e-3
rj2144 n949__vss n561__vss 114.4e-3
rj2145 n561__vss n656__vss 83.33e-3
rj2146 n949__vss n542__vss 114.4e-3
rj2147 n542__vss n657__vss 83.33e-3
rj2148 n949__vss n951__vss 103.3e-3
rj2149 n951__vss n529__vss 95.53e-3
rj2151 n951__vss n953__vss 65.33e-3
rj2152 n953__vss n516__vss 95.53e-3
rj2153 n516__vss n659__vss 83.33e-3
rj2154 n953__vss n954__vss 106.3e-3
rj2156 n954__vss n507__vss 114.4e-3
rj2158 n954__vss n490__vss 114.4e-3
rj2159 n490__vss n661__vss 83.33e-3
rj2160 n954__vss n957__vss 102.3e-3
rj2161 n957__vss n481__vss 95.53e-3
rj2163 n957__vss n959__vss 65.33e-3
rj2164 n959__vss n464__vss 95.53e-3
rj2165 n464__vss n663__vss 83.33e-3
rj2166 n959__vss n960__vss 107.3e-3
rj2168 n960__vss n451__vss 114.4e-3
rj2169 n451__vss n664__vss 83.33e-3
rj2170 n960__vss n442__vss 114.4e-3
rj2172 n960__vss n963__vss 103.3e-3
rj2173 n963__vss n425__vss 95.53e-3
rj2174 n425__vss n666__vss 83.33e-3
rj2175 n963__vss n964__vss 70.34e-3
rj2176 n964__vss n412__vss 95.53e-3
rj2178 n964__vss n966__vss 101.3e-3
rj2180 n966__vss n399__vss 114.4e-3
rj2181 n399__vss n668__vss 83.33e-3
rj2182 n966__vss n390__vss 114.4e-3
rj2183 n390__vss n669__vss 83.33e-3
rj2184 n966__vss n968__vss 102.3e-3
rj2185 n968__vss n377__vss 95.53e-3
rj2186 n377__vss n670__vss 83.33e-3
rj2187 n968__vss n969__vss 70.34e-3
rj2188 n969__vss n360__vss 95.53e-3
rj2190 n969__vss n971__vss 102.3e-3
rj2192 n971__vss n351__vss 114.4e-3
rj2194 n971__vss n338__vss 114.4e-3
rj2196 n971__vss n975__vss 101.3e-3
rj2197 n975__vss n325__vss 95.53e-3
rj2198 n325__vss n674__vss 83.33e-3
rj2199 n975__vss n976__vss 70.34e-3
rj2200 n976__vss n312__vss 95.53e-3
rj2202 n976__vss n978__vss 103.3e-3
rj2204 n978__vss n297__vss 114.4e-3
rj2206 n978__vss n282__vss 114.4e-3
rj2208 n978__vss n982__vss 100.3e-3
rj2209 n982__vss n269__vss 95.53e-3
rj2211 n982__vss n984__vss 70.34e-3
rj2212 n984__vss n260__vss 95.53e-3
rj2214 n984__vss n986__vss 104.3e-3
rj2216 n986__vss n247__vss 114.4e-3
rj2217 n247__vss n680__vss 83.33e-3
rj2218 n986__vss n234__vss 114.4e-3
rj2219 n234__vss n681__vss 83.33e-3
rj2220 n986__vss n988__vss 108.3e-3
rj2221 n988__vss n221__vss 95.53e-3
rj2223 n988__vss n990__vss 65.33e-3
rj2224 n990__vss n208__vss 95.53e-3
rj2225 n208__vss n683__vss 83.33e-3
rj2226 n990__vss n991__vss 101.3e-3
rj2228 n991__vss n191__vss 114.4e-3
rj2230 n991__vss n182__vss 114.4e-3
rj2231 n182__vss n685__vss 83.33e-3
rj2232 n991__vss n994__vss 107.3e-3
rj2233 n994__vss n165__vss 95.53e-3
rj2235 n994__vss n996__vss 65.33e-3
rj2236 n996__vss n152__vss 95.53e-3
rj2237 n152__vss n687__vss 83.33e-3
rj2238 n996__vss n997__vss 102.3e-3
rj2240 n997__vss n143__vss 114.4e-3
rj2242 n997__vss n126__vss 114.4e-3
rj2244 n997__vss n1001__vss 106.3e-3
rj2245 n1001__vss n113__vss 95.53e-3
rj2247 n1001__vss n1003__vss 65.33e-3
rj2248 n1003__vss n100__vss 95.53e-3
rj2249 n100__vss n691__vss 83.33e-3
rj2250 n1003__vss n1004__vss 103.3e-3
rj2252 n1004__vss n87__vss 114.4e-3
rj2254 n1004__vss n74__vss 114.4e-3
rj2255 n74__vss n693__vss 83.33e-3
rj2256 n1004__vss n1007__vss 105.3e-3
rj2257 n1007__vss n61__vss 95.53e-3
rj2259 n1007__vss n1009__vss 66.33e-3
rj2260 n1009__vss n48__vss 95.53e-3
rj2261 n48__vss n695__vss 83.33e-3
rj2262 n1009__vss n1010__vss 103.3e-3
rj2264 n1010__vss n35__vss 114.4e-3
rj2265 n35__vss n696__vss 83.33e-3
rj2266 n1010__vss n22__vss 114.4e-3
rj2268 n1010__vss n9__vss 202e-3
rj2270 n894__vss n884__vss 83.33e-3
rj2271 n896__vss n854__vss 83.33e-3
rj2272 n898__vss n828__vss 83.33e-3
rj2273 n899__vss n815__vss 83.33e-3
rj2274 n902__vss n776__vss 83.33e-3
rj2275 n903__vss n763__vss 83.33e-3
rj2276 n904__vss n754__vss 83.33e-3
rj2277 n905__vss n737__vss 83.33e-3
rj2278 n651__vss n626__vss 83.33e-3
rj2279 n652__vss n613__vss 83.33e-3
rj2280 n658__vss n529__vss 83.33e-3
rj2281 n660__vss n507__vss 83.33e-3
rj2282 n662__vss n481__vss 83.33e-3
rj2283 n665__vss n442__vss 83.33e-3
rj2284 n667__vss n412__vss 83.33e-3
rj2285 n671__vss n360__vss 83.33e-3
rj2286 n672__vss n351__vss 83.33e-3
rj2287 n673__vss n338__vss 83.33e-3
rj2288 n675__vss n312__vss 83.33e-3
rj2289 n676__vss n297__vss 83.33e-3
rj2290 n677__vss n282__vss 83.33e-3
rj2291 n678__vss n269__vss 83.33e-3
rj2292 n679__vss n260__vss 83.33e-3
rj2293 n682__vss n221__vss 83.33e-3
rj2294 n684__vss n191__vss 83.33e-3
rj2295 n686__vss n165__vss 83.33e-3
rj2296 n688__vss n143__vss 83.33e-3
rj2297 n689__vss n126__vss 83.33e-3
rj2298 n690__vss n113__vss 83.33e-3
rj2299 n692__vss n87__vss 83.33e-3
rj2300 n694__vss n61__vss 83.33e-3
rj2301 n697__vss n22__vss 83.33e-3
rj2303 n1507__vddio n1529__vddio 150.9e-3
rj2305 n1529__vddio n1531__vddio 90.27e-3
rj2306 n1531__vddio n1532__vddio 65.33e-3
rj2307 n1532__vddio n1533__vddio 49.2e-3
rj2309 n1533__vddio n1535__vddio 86.26e-3
rj2310 n1535__vddio n1536__vddio 70.34e-3
rj2311 n1536__vddio n1537__vddio 65.33e-3
rj2312 n1537__vddio n1538__vddio 50.2e-3
rj2314 n1538__vddio n1540__vddio 85.26e-3
rj2315 n1540__vddio n1541__vddio 70.34e-3
rj2316 n1541__vddio n1542__vddio 65.33e-3
rj2317 n1542__vddio n1543__vddio 51.2e-3
rj2319 n1543__vddio n1545__vddio 84.26e-3
rj2320 n1545__vddio n1546__vddio 70.34e-3
rj2321 n1546__vddio n1547__vddio 120.3e-3
rj2323 n1547__vddio n1549__vddio 105.3e-3
rj2324 n1549__vddio n1550__vddio 65.33e-3
rj2325 n1550__vddio n1551__vddio 104.3e-3
rj2327 n1551__vddio n1553__vddio 104.3e-3
rj2328 n1553__vddio n1554__vddio 65.33e-3
rj2329 n1554__vddio n1555__vddio 105.3e-3
rj2331 n1555__vddio n1557__vddio 103.3e-3
rj2332 n1557__vddio n1558__vddio 65.33e-3
rj2333 n1558__vddio n1559__vddio 106.3e-3
rj2335 n1559__vddio n1561__vddio 102.3e-3
rj2336 n1561__vddio n1562__vddio 65.33e-3
rj2337 n1562__vddio n1563__vddio 107.3e-3
rj2339 n1563__vddio n1565__vddio 103.3e-3
rj2340 n1565__vddio n1566__vddio 70.34e-3
rj2341 n1566__vddio n1567__vddio 101.3e-3
rj2343 n1567__vddio n1569__vddio 102.3e-3
rj2344 n1569__vddio n1570__vddio 70.34e-3
rj2345 n1570__vddio n1571__vddio 102.3e-3
rj2347 n1571__vddio n1573__vddio 101.3e-3
rj2348 n1573__vddio n1574__vddio 70.34e-3
rj2349 n1574__vddio n1575__vddio 103.3e-3
rj2351 n1575__vddio n1577__vddio 100.3e-3
rj2352 n1577__vddio n1578__vddio 70.34e-3
rj2353 n1578__vddio n1579__vddio 104.3e-3
rj2355 n1579__vddio n1581__vddio 108.3e-3
rj2356 n1581__vddio n1582__vddio 65.33e-3
rj2357 n1582__vddio n1583__vddio 101.3e-3
rj2359 n1583__vddio n1585__vddio 107.3e-3
rj2360 n1585__vddio n1586__vddio 65.33e-3
rj2361 n1586__vddio n1587__vddio 102.3e-3
rj2363 n1587__vddio n1589__vddio 106.3e-3
rj2364 n1589__vddio n1590__vddio 65.33e-3
rj2365 n1590__vddio n1591__vddio 103.3e-3
rj2367 n1591__vddio n1593__vddio 105.3e-3
rj2368 n1593__vddio n1594__vddio 66.33e-3
rj2369 n1594__vddio n1595__vddio 103.3e-3
rj2371 n1595__vddio n14__vddio 205.7e-3
rj2373 n1529__vddio n1492__vddio 118.1e-3
rj2375 n1531__vddio n1464__vddio 99.2e-3
rj2376 n1464__vddio n1509__vddio 83.33e-3
rj2377 n1532__vddio n1443__vddio 99.2e-3
rj2379 n1533__vddio n1422__vddio 118.1e-3
rj2380 n1422__vddio n1511__vddio 83.33e-3
rj2381 n1535__vddio n1391__vddio 99.2e-3
rj2383 n1536__vddio n1370__vddio 99.2e-3
rj2385 n1537__vddio n1356__vddio 99.2e-3
rj2386 n1356__vddio n1514__vddio 83.33e-3
rj2387 n1538__vddio n1328__vddio 118.1e-3
rj2388 n1328__vddio n1515__vddio 83.33e-3
rj2389 n1540__vddio n1307__vddio 99.2e-3
rj2391 n1541__vddio n1276__vddio 99.2e-3
rj2393 n1542__vddio n1262__vddio 99.2e-3
rj2395 n1543__vddio n1234__vddio 118.1e-3
rj2397 n1545__vddio n1213__vddio 99.2e-3
rj2398 n1213__vddio n1520__vddio 83.33e-3
rj2399 n1546__vddio n1186__vddio 99.2e-3
rj2401 n1549__vddio n1112__vddio 99.2e-3
rj2403 n1550__vddio n1091__vddio 99.2e-3
rj2405 n1551__vddio n1070__vddio 118.1e-3
rj2406 n1070__vddio n1122__vddio 83.33e-3
rj2407 n1551__vddio n1049__vddio 118.1e-3
rj2409 n1553__vddio n1025__vddio 99.2e-3
rj2410 n1025__vddio n1124__vddio 83.33e-3
rj2411 n1554__vddio n997__vddio 99.2e-3
rj2412 n997__vddio n1125__vddio 83.33e-3
rj2413 n1555__vddio n976__vddio 118.1e-3
rj2415 n1555__vddio n955__vddio 118.1e-3
rj2417 n1557__vddio n934__vddio 99.2e-3
rj2419 n1558__vddio n903__vddio 99.2e-3
rj2420 n903__vddio n1129__vddio 83.33e-3
rj2421 n1559__vddio n889__vddio 118.1e-3
rj2423 n1559__vddio n861__vddio 118.1e-3
rj2424 n861__vddio n1131__vddio 83.33e-3
rj2425 n1561__vddio n847__vddio 99.2e-3
rj2427 n1562__vddio n813__vddio 99.2e-3
rj2428 n813__vddio n1133__vddio 83.33e-3
rj2429 n1563__vddio n788__vddio 118.1e-3
rj2430 n788__vddio n1134__vddio 83.33e-3
rj2431 n1563__vddio n767__vddio 118.1e-3
rj2433 n1565__vddio n746__vddio 99.2e-3
rj2434 n746__vddio n1136__vddio 83.33e-3
rj2435 n1566__vddio n725__vddio 99.2e-3
rj2437 n1567__vddio n704__vddio 118.1e-3
rj2438 n704__vddio n1138__vddio 83.33e-3
rj2439 n1567__vddio n690__vddio 118.1e-3
rj2440 n690__vddio n1139__vddio 83.33e-3
rj2441 n1569__vddio n662__vddio 99.2e-3
rj2442 n662__vddio n1140__vddio 83.33e-3
rj2443 n1570__vddio n631__vddio 99.2e-3
rj2445 n1571__vddio n617__vddio 118.1e-3
rj2447 n1571__vddio n589__vddio 118.1e-3
rj2449 n1573__vddio n565__vddio 99.2e-3
rj2450 n565__vddio n1144__vddio 83.33e-3
rj2451 n1574__vddio n537__vddio 99.2e-3
rj2453 n1575__vddio n516__vddio 118.1e-3
rj2455 n1575__vddio n495__vddio 118.1e-3
rj2457 n1577__vddio n474__vddio 99.2e-3
rj2459 n1578__vddio n454__vddio 99.2e-3
rj2461 n1579__vddio n433__vddio 118.1e-3
rj2462 n433__vddio n1150__vddio 83.33e-3
rj2463 n1579__vddio n408__vddio 118.1e-3
rj2465 n1581__vddio n387__vddio 99.2e-3
rj2466 n387__vddio n1152__vddio 83.33e-3
rj2467 n1582__vddio n366__vddio 99.2e-3
rj2469 n1583__vddio n338__vddio 118.1e-3
rj2470 n338__vddio n1154__vddio 83.33e-3
rj2471 n1583__vddio n324__vddio 118.1e-3
rj2473 n1585__vddio n296__vddio 99.2e-3
rj2474 n296__vddio n1156__vddio 83.33e-3
rj2475 n1586__vddio n265__vddio 99.2e-3
rj2476 n265__vddio n1157__vddio 83.33e-3
rj2477 n1587__vddio n251__vddio 118.1e-3
rj2479 n1587__vddio n223__vddio 118.1e-3
rj2481 n1589__vddio n192__vddio 99.2e-3
rj2483 n1590__vddio n171__vddio 99.2e-3
rj2484 n171__vddio n1161__vddio 83.33e-3
rj2485 n1591__vddio n150__vddio 118.1e-3
rj2487 n1591__vddio n129__vddio 118.1e-3
rj2488 n129__vddio n1163__vddio 83.33e-3
rj2489 n1593__vddio n108__vddio 99.2e-3
rj2491 n1594__vddio n81__vddio 99.2e-3
rj2492 n81__vddio n1165__vddio 83.33e-3
rj2493 n1595__vddio n56__vddio 118.1e-3
rj2494 n56__vddio n1166__vddio 83.33e-3
rj2495 n1595__vddio n35__vddio 118.1e-3
rj2497 n1508__vddio n1492__vddio 83.33e-3
rj2498 n1510__vddio n1443__vddio 83.33e-3
rj2499 n1512__vddio n1391__vddio 83.33e-3
rj2500 n1513__vddio n1370__vddio 83.33e-3
rj2501 n1516__vddio n1307__vddio 83.33e-3
rj2502 n1517__vddio n1276__vddio 83.33e-3
rj2503 n1518__vddio n1262__vddio 83.33e-3
rj2504 n1519__vddio n1234__vddio 83.33e-3
rj2505 n1121__vddio n1091__vddio 83.33e-3
rj2506 n1123__vddio n1049__vddio 83.33e-3
rj2507 n1126__vddio n976__vddio 83.33e-3
rj2508 n1127__vddio n955__vddio 83.33e-3
rj2509 n1128__vddio n934__vddio 83.33e-3
rj2510 n1130__vddio n889__vddio 83.33e-3
rj2511 n1132__vddio n847__vddio 83.33e-3
rj2512 n1135__vddio n767__vddio 83.33e-3
rj2513 n1137__vddio n725__vddio 83.33e-3
rj2514 n1141__vddio n631__vddio 83.33e-3
rj2515 n1142__vddio n617__vddio 83.33e-3
rj2516 n1143__vddio n589__vddio 83.33e-3
rj2517 n1145__vddio n537__vddio 83.33e-3
rj2518 n1146__vddio n516__vddio 83.33e-3
rj2519 n1147__vddio n495__vddio 83.33e-3
rj2520 n1148__vddio n474__vddio 83.33e-3
rj2521 n1149__vddio n454__vddio 83.33e-3
rj2522 n1151__vddio n408__vddio 83.33e-3
rj2523 n1153__vddio n366__vddio 83.33e-3
rj2524 n1155__vddio n324__vddio 83.33e-3
rj2525 n1158__vddio n251__vddio 83.33e-3
rj2526 n1159__vddio n223__vddio 83.33e-3
rj2527 n1160__vddio n192__vddio 83.33e-3
rj2528 n1162__vddio n150__vddio 83.33e-3
rj2529 n1164__vddio n108__vddio 83.33e-3
rj2530 n1167__vddio n35__vddio 83.33e-3
rj2531 n61__i1__i13__net1 n63__i1__i13__net1 125e-3
rj2532 n64__i1__i13__net1 n62__i1__i13__net1 125e-3
rj2533 n29__i1__i12__net1 n31__i1__i12__net1 125e-3
rj2534 n32__i1__i12__net1 n30__i1__i12__net1 125e-3
rj2535 n8__i1__i13__net1 n63__i1__i13__net1 250e-3
rj2536 n64__i1__i13__net1 n6__i1__i13__net1 250e-3
rj2537 n33__i1__i12__net1 n35__i1__i12__net1 125e-3
rj2538 n36__i1__i12__net1 n34__i1__i12__net1 125e-3
rj2539 n75__i1__i13__net1 n73__i1__i13__net1 125e-3
rj2540 n74__i1__i13__net1 n76__i1__i13__net1 125e-3
rj2541 n39__i1__i12__net1 n37__i1__i12__net1 125e-3
rj2542 n38__i1__i12__net1 n40__i1__i12__net1 125e-3
rj2543 n75__i1__i13__net1 n85__i1__i13__net1 125e-3
rj2544 n86__i1__i13__net1 n76__i1__i13__net1 125e-3
rj2545 n43__i1__i12__net1 n41__i1__i12__net1 125e-3
rj2546 n42__i1__i12__net1 n44__i1__i12__net1 125e-3
rj2547 n93__i1__i13__net1 n20__i1__i13__net1 250e-3
rj2548 n18__i1__i13__net1 n96__i1__i13__net1 250e-3
rj2549 n43__i1__i12__net1 n45__i1__i12__net1 125e-3
rj2550 n46__i1__i12__net1 n44__i1__i12__net1 125e-3
rj2551 n101__i1__i13__net1 n93__i1__i13__net1 125e-3
rj2552 n96__i1__i13__net1 n102__i1__i13__net1 125e-3
rj2553 n49__i1__i12__net1 n51__i1__i12__net1 125e-3
rj2554 n52__i1__i12__net1 n50__i1__i12__net1 125e-3
rj2555 n105__i1__i13__net1 n27__i1__i13__net1 250e-3
rj2556 n26__i1__i13__net1 n108__i1__i13__net1 250e-3
rj2557 n51__i1__i12__net1 n26__i1__i12__net1 250e-3
rj2558 n28__i1__i12__net1 n52__i1__i12__net1 250e-3
rj2559 n105__i1__i13__net1 n32__i1__i13__net1 250e-3
rj2560 n30__i1__i13__net1 n108__i1__i13__net1 250e-3
rj2561 n113__i1__i13__net1 n115__i1__i13__net1 125e-3
rj2562 n116__i1__i13__net1 n114__i1__i13__net1 125e-3
rj2563 n117__i1__i13__net1 n115__i1__i13__net1 125e-3
rj2564 n116__i1__i13__net1 n118__i1__i13__net1 125e-3
rj2565 n15__i1__net4 n13__i1__net4 125e-3
rj2566 n14__i1__net4 n15__i1__net4 125e-3
rj2567 n65__i1__i12__net1 n57__i1__i12__net1 231e-3
rj2568 n57__i1__i12__net1 n64__i1__i12__net1 237.5e-3
rj2569 n127__i1__i13__net1 n125__i1__i13__net1 125e-3
rj2570 n126__i1__i13__net1 n128__i1__i13__net1 125e-3
rj2571 n17__i1__net4 n19__i1__net4 125e-3
rj2572 n19__i1__net4 n18__i1__net4 125e-3
rj2573 n129__i1__i13__net1 n127__i1__i13__net1 125e-3
rj2574 n128__i1__i13__net1 n130__i1__i13__net1 125e-3
rj2576 n1584__vss n1586__vss 330.5e-3
rj2577 n1586__vss n1577__vss 12.5e-3
rj2578 n1573__vss n1584__vss 25e-3
rj2580 n1730__vddio n1732__vddio 210.4e-3
rj2581 n1732__vddio n1733__vddio 8.333e-3
rj2582 n133__i1__i13__net1 n135__i1__i13__net1 125e-3
rj2583 n136__i1__i13__net1 n134__i1__i13__net1 125e-3
rj2584 n135__i1__i13__net1 n137__i1__i13__net1 125e-3
rj2585 n138__i1__i13__net1 n136__i1__i13__net1 125e-3
rj2586 n141__i1__i13__net1 n143__i1__i13__net1 125e-3
rj2587 n144__i1__i13__net1 n142__i1__i13__net1 125e-3
rj2588 n143__i1__i13__net1 n68__i1__i13__net1 250e-3
rj2589 n66__i1__i13__net1 n144__i1__i13__net1 250e-3
rj2590 n26__piso_out n31__piso_out 304.1e-3
rj2591 n31__piso_out n29__piso_out 33.55e-3
rj2592 n29__piso_out n28__piso_out 34.46e-3
rj2593 n149__i1__i13__net1 n192__i1__i13__net1 125e-3
rj2594 n193__i1__i13__net1 n150__i1__i13__net1 125e-3
rj2595 n192__i1__i13__net1 n151__i1__i13__net1 125e-3
rj2596 n152__i1__i13__net1 n193__i1__i13__net1 125e-3
rj2597 n196__i1__i13__net1 n153__i1__i13__net1 125e-3
rj2598 n154__i1__i13__net1 n197__i1__i13__net1 125e-3
rj2599 n155__i1__i13__net1 n196__i1__i13__net1 125e-3
rj2600 n197__i1__i13__net1 n156__i1__i13__net1 125e-3
rj2601 n23__i1__net4 n28__i1__net4 34e-3
rj2602 n28__i1__net4 n22__i1__net4 35.8e-3
rj2603 n22__i1__net4 n21__i1__net4 110.8e-3
rj2604 n28__i1__net4 n25__i1__net4 573.2e-3
rj2605 n229__i1__net2 n329__i1__net2 58.34e-3
rj2606 n329__i1__net2 n330__i1__net2 83.65e-3
rj2607 n330__i1__net2 n331__i1__net2 86.1e-3
rj2608 n331__i1__net2 n332__i1__net2 84.87e-3
rj2609 n332__i1__net2 n333__i1__net2 83.65e-3
rj2610 n333__i1__net2 n334__i1__net2 86.1e-3
rj2611 n334__i1__net2 n335__i1__net2 84.87e-3
rj2612 n335__i1__net2 n336__i1__net2 83.65e-3
rj2613 n336__i1__net2 n337__i1__net2 84.87e-3
rj2614 n337__i1__net2 n338__i1__net2 84.87e-3
rj2615 n338__i1__net2 n321__i1__net2 167e-3
rj2616 n236__i1__net2 n329__i1__net2 83.33e-3
rj2617 n240__i1__net2 n330__i1__net2 83.33e-3
rj2618 n254__i1__net2 n331__i1__net2 83.33e-3
rj2619 n263__i1__net2 n332__i1__net2 83.33e-3
rj2620 n272__i1__net2 n333__i1__net2 83.33e-3
rj2621 n281__i1__net2 n334__i1__net2 83.33e-3
rj2622 n290__i1__net2 n335__i1__net2 83.33e-3
rj2623 n299__i1__net2 n336__i1__net2 83.33e-3
rj2624 n308__i1__net2 n337__i1__net2 83.33e-3
rj2625 n312__i1__net2 n338__i1__net2 83.33e-3
rj2626 n228__i1__net2 n238__i1__net2 120.8e-3
rj2627 n238__i1__net2 n242__i1__net2 83.65e-3
rj2628 n242__i1__net2 n256__i1__net2 86.1e-3
rj2629 n256__i1__net2 n265__i1__net2 84.87e-3
rj2630 n265__i1__net2 n274__i1__net2 83.65e-3
rj2631 n274__i1__net2 n283__i1__net2 86.1e-3
rj2632 n283__i1__net2 n292__i1__net2 84.87e-3
rj2633 n292__i1__net2 n301__i1__net2 83.65e-3
rj2634 n301__i1__net2 n310__i1__net2 84.87e-3
rj2635 n310__i1__net2 n314__i1__net2 84.87e-3
rj2636 n314__i1__net2 n323__i1__net2 83.65e-3
rj2637 n15__piso_outinv n16__piso_outinv 70.81e-3
rj2638 n16__piso_outinv n18__piso_outinv 3.873e-3
rj2639 n18__piso_outinv n17__piso_outinv 47.35e-3
rj2640 n227__i1__net2 n339__i1__net2 120.8e-3
rj2641 n339__i1__net2 n340__i1__net2 86.1e-3
rj2642 n340__i1__net2 n341__i1__net2 83.65e-3
rj2643 n341__i1__net2 n342__i1__net2 84.87e-3
rj2644 n342__i1__net2 n343__i1__net2 83.65e-3
rj2645 n343__i1__net2 n344__i1__net2 86.1e-3
rj2646 n344__i1__net2 n345__i1__net2 84.87e-3
rj2647 n345__i1__net2 n346__i1__net2 83.65e-3
rj2648 n346__i1__net2 n347__i1__net2 84.87e-3
rj2649 n347__i1__net2 n348__i1__net2 86.1e-3
rj2650 n348__i1__net2 n324__i1__net2 168.2e-3
rj2651 n230__i1__net2 n339__i1__net2 83.33e-3
rj2652 n243__i1__net2 n340__i1__net2 83.33e-3
rj2653 n248__i1__net2 n341__i1__net2 83.33e-3
rj2654 n257__i1__net2 n342__i1__net2 83.33e-3
rj2655 n266__i1__net2 n343__i1__net2 83.33e-3
rj2656 n275__i1__net2 n344__i1__net2 83.33e-3
rj2657 n284__i1__net2 n345__i1__net2 83.33e-3
rj2658 n293__i1__net2 n346__i1__net2 83.33e-3
rj2659 n302__i1__net2 n347__i1__net2 83.33e-3
rj2660 n315__i1__net2 n348__i1__net2 83.33e-3
rj2661 n226__i1__net2 n349__i1__net2 120.8e-3
rj2662 n349__i1__net2 n350__i1__net2 86.1e-3
rj2663 n350__i1__net2 n351__i1__net2 83.65e-3
rj2664 n351__i1__net2 n352__i1__net2 84.87e-3
rj2665 n352__i1__net2 n353__i1__net2 83.65e-3
rj2666 n353__i1__net2 n354__i1__net2 86.1e-3
rj2667 n354__i1__net2 n355__i1__net2 84.87e-3
rj2668 n355__i1__net2 n356__i1__net2 83.65e-3
rj2669 n356__i1__net2 n357__i1__net2 84.87e-3
rj2670 n357__i1__net2 n358__i1__net2 86.1e-3
rj2671 n358__i1__net2 n325__i1__net2 168.2e-3
rj2672 n231__i1__net2 n349__i1__net2 83.33e-3
rj2673 n244__i1__net2 n350__i1__net2 83.33e-3
rj2674 n249__i1__net2 n351__i1__net2 83.33e-3
rj2675 n258__i1__net2 n352__i1__net2 83.33e-3
rj2676 n267__i1__net2 n353__i1__net2 83.33e-3
rj2677 n276__i1__net2 n354__i1__net2 83.33e-3
rj2678 n285__i1__net2 n355__i1__net2 83.33e-3
rj2679 n294__i1__net2 n356__i1__net2 83.33e-3
rj2680 n303__i1__net2 n357__i1__net2 83.33e-3
rj2681 n316__i1__net2 n358__i1__net2 83.33e-3
rj2682 n225__i1__net2 n234__i1__net2 120.8e-3
rj2683 n234__i1__net2 n247__i1__net2 86.1e-3
rj2684 n247__i1__net2 n252__i1__net2 83.65e-3
rj2685 n252__i1__net2 n261__i1__net2 84.87e-3
rj2686 n261__i1__net2 n270__i1__net2 83.65e-3
rj2687 n270__i1__net2 n279__i1__net2 86.1e-3
rj2688 n279__i1__net2 n288__i1__net2 84.87e-3
rj2689 n288__i1__net2 n297__i1__net2 83.65e-3
rj2690 n297__i1__net2 n306__i1__net2 84.87e-3
rj2691 n306__i1__net2 n319__i1__net2 86.1e-3
rj2692 n319__i1__net2 n328__i1__net2 84.87e-3
rj2693 n200__i1__i13__net1 n157__i1__i13__net1 125e-3
rj2694 n158__i1__i13__net1 n201__i1__i13__net1 125e-3
rj2696 n1664__vss n1666__vss 550.8e-3
rj2697 n1666__vss n1617__vss 25e-3
rj2698 n1614__vss n1664__vss 500e-3
rj2699 n7__i1__i11__outinv n11__i1__i11__outinv 1.0562
rj2700 n11__i1__i11__outinv n10__i1__i11__outinv 92.37e-3
rj2701 n66__i1__net3 n54__i1__net3 125e-3
rj2702 n55__i1__net3 n67__i1__net3 125e-3
rj2703 n66__i1__net3 n56__i1__net3 125e-3
rj2704 n57__i1__net3 n67__i1__net3 125e-3
rj2705 n70__i1__net3 n58__i1__net3 125e-3
rj2706 n59__i1__net3 n70__i1__net3 125e-3
rj2707 n72__i1__net3 n60__i1__net3 125e-3
rj2708 n61__i1__net3 n72__i1__net3 125e-3
rj2709 n74__i1__net3 n62__i1__net3 125e-3
rj2710 n63__i1__net3 n74__i1__net3 125e-3
rj2711 n202__i1__i13__net1 n203__i1__i13__net1 156.3e-3
rj2712 n203__i1__i13__net1 n204__i1__i13__net1 86.1e-3
rj2713 n204__i1__i13__net1 n182__i1__i13__net1 168.2e-3
rj2714 n160__i1__i13__net1 n203__i1__i13__net1 83.33e-3
rj2715 n171__i1__i13__net1 n204__i1__i13__net1 83.33e-3
rj2716 n205__i1__i13__net1 n162__i1__i13__net1 156.3e-3
rj2717 n162__i1__i13__net1 n173__i1__i13__net1 86.1e-3
rj2718 n173__i1__i13__net1 n184__i1__i13__net1 84.87e-3
rj2719 n206__i1__i13__net1 n207__i1__i13__net1 156.3e-3
rj2720 n207__i1__i13__net1 n208__i1__i13__net1 86.1e-3
rj2721 n208__i1__i13__net1 n190__i1__i13__net1 168.2e-3
rj2722 n168__i1__i13__net1 n207__i1__i13__net1 83.33e-3
rj2723 n179__i1__i13__net1 n208__i1__i13__net1 83.33e-3
rj2724 n209__i1__i13__net1 n210__i1__i13__net1 155.1e-3
rj2725 n210__i1__i13__net1 n211__i1__i13__net1 86.1e-3
rj2726 n211__i1__i13__net1 n189__i1__i13__net1 168.2e-3
rj2727 n167__i1__i13__net1 n210__i1__i13__net1 83.33e-3
rj2728 n178__i1__i13__net1 n211__i1__i13__net1 83.33e-3
rj2729 n212__i1__i13__net1 n213__i1__i13__net1 155.1e-3
rj2730 n213__i1__i13__net1 n214__i1__i13__net1 86.1e-3
rj2731 n214__i1__i13__net1 n186__i1__i13__net1 168.2e-3
rj2732 n164__i1__i13__net1 n213__i1__i13__net1 83.33e-3
rj2733 n175__i1__i13__net1 n214__i1__i13__net1 83.33e-3
rj2734 n76__i1__net3 n64__i1__net3 125e-3
rj2735 n65__i1__net3 n76__i1__net3 125e-3
rj2737 n1656__vss n1647__vss 114.9e-3
rj2739 n1647__vss n1669__vss 110e-3
rj2741 n1669__vss n1637__vss 114.9e-3
rj2743 n1637__vss n1672__vss 178.3e-3
rj2745 n1672__vss n1612__vss 114.9e-3
rj2747 n1612__vss n1675__vss 110e-3
rj2749 n1675__vss n1600__vss 114.9e-3
rj2751 n1600__vss n1678__vss 111.6e-3
rj2753 n1678__vss n1570__vss 114.9e-3
rj2755 n1570__vss n1681__vss 110e-3
rj2757 n1681__vss n1559__vss 114.9e-3
rj2759 n1559__vss n1310__vss 114.9e-3
rj2761 n1310__vss n1303__vss 114.9e-3
rj2763 n1303__vss n1686__vss 110e-3
rj2764 n1686__vss n1687__vss 125e-3
rj2765 n1641__vss n1669__vss 125e-3
rj2766 n1624__vss n1672__vss 125e-3
rj2767 n1604__vss n1675__vss 125e-3
rj2768 n1587__vss n1678__vss 125e-3
rj2769 n1563__vss n1681__vss 125e-3
rj2770 n1292__vss n1686__vss 125e-3
rj2772 n1813__vddio n1828__vddio 114.9e-3
rj2774 n1828__vddio n1830__vddio 110e-3
rj2776 n1830__vddio n1792__vddio 114.9e-3
rj2778 n1792__vddio n1833__vddio 178.3e-3
rj2780 n1833__vddio n1835__vddio 114.9e-3
rj2782 n1835__vddio n1837__vddio 110e-3
rj2784 n1837__vddio n1839__vddio 114.9e-3
rj2786 n1839__vddio n1841__vddio 111.6e-3
rj2788 n1841__vddio n1843__vddio 114.9e-3
rj2790 n1843__vddio n1706__vddio 110e-3
rj2792 n1706__vddio n1846__vddio 115.4e-3
rj2794 n1846__vddio n1848__vddio 115.4e-3
rj2796 n1848__vddio n1850__vddio 112.2e-3
rj2798 n1850__vddio n1852__vddio 113.8e-3
rj2799 n1852__vddio n1684__vddio 125e-3
rj2800 n1812__vddio n1828__vddio 125e-3
rj2801 n1805__vddio n1830__vddio 125e-3
rj2802 n1791__vddio n1833__vddio 125e-3
rj2803 n1765__vddio n1835__vddio 125e-3
rj2804 n1758__vddio n1837__vddio 125e-3
rj2805 n1751__vddio n1839__vddio 125e-3
rj2806 n1744__vddio n1841__vddio 125e-3
rj2807 n1719__vddio n1843__vddio 125e-3
rj2808 n1705__vddio n1846__vddio 125e-3
rj2809 n1698__vddio n1848__vddio 125e-3
rj2810 n1691__vddio n1850__vddio 125e-3
rj2811 n1652__vss n1688__vss 168.2e-3
rj2812 n1688__vss n1689__vss 86.1e-3
rj2813 n1689__vss n1690__vss 84.87e-3
rj2814 n1690__vss n1691__vss 130.1e-3
rj2815 n1691__vss n1692__vss 87.32e-3
rj2816 n1692__vss n1693__vss 83.65e-3
rj2817 n1693__vss n1694__vss 84.87e-3
rj2818 n1694__vss n1695__vss 83.65e-3
rj2819 n1695__vss n1696__vss 84.87e-3
rj2820 n1696__vss n1697__vss 86.1e-3
rj2821 n1697__vss n1698__vss 83.65e-3
rj2822 n1698__vss n1699__vss 84.87e-3
rj2823 n1699__vss n1700__vss 84.87e-3
rj2824 n1700__vss n1295__vss 168.2e-3
rj2825 n1644__vss n1688__vss 83.33e-3
rj2826 n1638__vss n1689__vss 83.33e-3
rj2827 n1633__vss n1690__vss 83.33e-3
rj2828 n1627__vss n1691__vss 83.33e-3
rj2829 n1610__vss n1692__vss 83.33e-3
rj2830 n1601__vss n1693__vss 83.33e-3
rj2831 n1596__vss n1694__vss 83.33e-3
rj2832 n1590__vss n1695__vss 83.33e-3
rj2833 n1566__vss n1696__vss 83.33e-3
rj2834 n1560__vss n1697__vss 83.33e-3
rj2835 n1555__vss n1698__vss 83.33e-3
rj2836 n1306__vss n1699__vss 83.33e-3
rj2837 n1299__vss n1700__vss 83.33e-3
rj2838 n1654__vss n1649__vss 168.2e-3
rj2839 n1649__vss n1643__vss 86.1e-3
rj2840 n1643__vss n1701__vss 84.87e-3
rj2841 n1701__vss n1702__vss 130.1e-3
rj2842 n1702__vss n1607__vss 86.1e-3
rj2843 n1607__vss n1606__vss 84.87e-3
rj2844 n1606__vss n1703__vss 84.87e-3
rj2845 n1703__vss n1704__vss 83.65e-3
rj2846 n1704__vss n1571__vss 84.87e-3
rj2847 n1571__vss n1565__vss 86.1e-3
rj2848 n1565__vss n1705__vss 83.65e-3
rj2849 n1705__vss n1311__vss 84.87e-3
rj2850 n1311__vss n1304__vss 86.1e-3
rj2851 n1304__vss n1297__vss 167e-3
rj2852 n1635__vss n1701__vss 83.33e-3
rj2853 n1629__vss n1702__vss 83.33e-3
rj2854 n1598__vss n1703__vss 83.33e-3
rj2855 n1592__vss n1704__vss 83.33e-3
rj2856 n1557__vss n1705__vss 83.33e-3
rj2857 n1819__vddio n1806__vddio 84.87e-3
rj2858 n1806__vddio n1799__vddio 86.1e-3
rj2859 n1799__vddio n1798__vddio 84.87e-3
rj2860 n1798__vddio n1785__vddio 130.1e-3
rj2861 n1785__vddio n1759__vddio 84.87e-3
rj2862 n1759__vddio n1752__vddio 86.1e-3
rj2863 n1752__vddio n1745__vddio 84.87e-3
rj2864 n1745__vddio n1738__vddio 83.65e-3
rj2865 n1738__vddio n1713__vddio 84.87e-3
rj2866 n1713__vddio n1712__vddio 86.1e-3
rj2867 n1712__vddio n1699__vddio 83.65e-3
rj2868 n1699__vddio n1692__vddio 84.87e-3
rj2869 n1692__vddio n1685__vddio 83.65e-3
rj2870 n1685__vddio n1678__vddio 86.1e-3
rj2871 n1817__vddio n1853__vddio 168.2e-3
rj2872 n1853__vddio n1854__vddio 86.1e-3
rj2873 n1854__vddio n1855__vddio 84.87e-3
rj2874 n1855__vddio n1856__vddio 130.1e-3
rj2875 n1856__vddio n1857__vddio 84.87e-3
rj2876 n1857__vddio n1858__vddio 86.1e-3
rj2877 n1858__vddio n1859__vddio 84.87e-3
rj2878 n1859__vddio n1860__vddio 83.65e-3
rj2879 n1860__vddio n1861__vddio 84.87e-3
rj2880 n1861__vddio n1862__vddio 86.1e-3
rj2881 n1862__vddio n1863__vddio 83.65e-3
rj2882 n1863__vddio n1864__vddio 84.87e-3
rj2883 n1864__vddio n1865__vddio 83.65e-3
rj2884 n1865__vddio n1681__vddio 169.4e-3
rj2885 n1809__vddio n1853__vddio 83.33e-3
rj2886 n1802__vddio n1854__vddio 83.33e-3
rj2887 n1796__vddio n1855__vddio 83.33e-3
rj2888 n1788__vddio n1856__vddio 83.33e-3
rj2889 n1762__vddio n1857__vddio 83.33e-3
rj2890 n1755__vddio n1858__vddio 83.33e-3
rj2891 n1748__vddio n1859__vddio 83.33e-3
rj2892 n1741__vddio n1860__vddio 83.33e-3
rj2893 n1716__vddio n1861__vddio 83.33e-3
rj2894 n1710__vddio n1862__vddio 83.33e-3
rj2895 n1702__vddio n1863__vddio 83.33e-3
rj2896 n1695__vddio n1864__vddio 83.33e-3
rj2897 n1688__vddio n1865__vddio 83.33e-3
rj2898 n1814__vddio n1866__vddio 168.2e-3
rj2899 n1866__vddio n1867__vddio 86.1e-3
rj2900 n1867__vddio n1868__vddio 84.87e-3
rj2901 n1868__vddio n1869__vddio 130.1e-3
rj2902 n1869__vddio n1870__vddio 84.87e-3
rj2903 n1870__vddio n1871__vddio 86.1e-3
rj2904 n1871__vddio n1872__vddio 84.87e-3
rj2905 n1872__vddio n1873__vddio 83.65e-3
rj2906 n1873__vddio n1874__vddio 84.87e-3
rj2907 n1874__vddio n1875__vddio 86.1e-3
rj2908 n1875__vddio n1876__vddio 83.65e-3
rj2909 n1876__vddio n1877__vddio 84.87e-3
rj2910 n1877__vddio n1878__vddio 83.65e-3
rj2911 n1878__vddio n1683__vddio 169.4e-3
rj2912 n1811__vddio n1866__vddio 83.33e-3
rj2913 n1804__vddio n1867__vddio 83.33e-3
rj2914 n1793__vddio n1868__vddio 83.33e-3
rj2915 n1790__vddio n1869__vddio 83.33e-3
rj2916 n1764__vddio n1870__vddio 83.33e-3
rj2917 n1757__vddio n1871__vddio 83.33e-3
rj2918 n1750__vddio n1872__vddio 83.33e-3
rj2919 n1743__vddio n1873__vddio 83.33e-3
rj2920 n1718__vddio n1874__vddio 83.33e-3
rj2921 n1707__vddio n1875__vddio 83.33e-3
rj2922 n1704__vddio n1876__vddio 83.33e-3
rj2923 n1697__vddio n1877__vddio 83.33e-3
rj2924 n1690__vddio n1878__vddio 83.33e-3
rj2926 n1879__vddio n1881__vddio 259.5e-3
rj2928 n1881__vddio n1883__vddio 280.5e-3
rj2930 n1883__vddio n1885__vddio 280.5e-3
rj2931 n1885__vddio n1826__vddio 8.333e-3
rj2932 n1820__vddio n1879__vddio 9.804e-3
rj2933 n1822__vddio n1881__vddio 8.333e-3
rj2934 n1824__vddio n1883__vddio 8.333e-3
rj2936 n1706__vss n1708__vss 259.5e-3
rj2938 n1708__vss n1710__vss 280.5e-3
rj2940 n1710__vss n1712__vss 280.5e-3
rj2941 n1712__vss n1713__vss 8.333e-3
rj2942 n1657__vss n1706__vss 9.804e-3
rj2943 n1659__vss n1708__vss 8.333e-3
rj2944 n1661__vss n1710__vss 8.333e-3
rj2945 n1663__vss n1712__vss 8.333e-3
rj2946 n78__i1__net3 n79__i1__net3 1.7714
rj2947 n79__i1__net3 n80__i1__net3 38.53e-3
rj2948 n79__i1__net3 i1__net3 205.1e-3
rj2949 i1__net3 n81__i1__net3 110.6e-3
rj2950 n81__i1__net3 n17__i1__net3 113.8e-3
rj2951 n17__i1__net3 n28__i1__net3 115.4e-3
rj2952 n80__i1__net3 n82__i1__net3 110.6e-3
rj2953 n82__i1__net3 n83__i1__net3 114.9e-3
rj2954 n83__i1__net3 n26__i1__net3 236.6e-3
rj2955 n6__i1__net3 n80__i1__net3 125e-3
rj2956 n8__i1__net3 n81__i1__net3 125e-3
rj2957 n14__i1__net3 n82__i1__net3 125e-3
rj2958 n21__i1__net3 n83__i1__net3 125e-3
rk2 n2__chipdriverout n4__chipdriverout 126.2e-3
rk3 n4__chipdriverout n5__chipdriverout 237.9e-3
rk4 n5__chipdriverout n6__chipdriverout 344.7e-3
rk5 n6__chipdriverout n7__chipdriverout 142.4e-3
rk6 n7__chipdriverout n8__chipdriverout 225e-3
rk7 n8__chipdriverout n9__chipdriverout 360.9e-3
rk8 n9__chipdriverout n10__chipdriverout 139.1e-3
rk9 n10__chipdriverout n11__chipdriverout 226.6e-3
rk10 n11__chipdriverout n12__chipdriverout 341.4e-3
rk11 n12__chipdriverout n13__chipdriverout 157e-3
rk12 n13__chipdriverout n14__chipdriverout 303.3e-3
rk13 n3__chipdriverout n4__chipdriverout 3.1
rk14 n3__chipdriverout n7__chipdriverout 3.1
rk15 n3__chipdriverout n10__chipdriverout 3.1
rk16 n3__chipdriverout n13__chipdriverout 3.1
rk18 n17__chipdriverout n18__chipdriverout 10.04e-3
rk19 n18__chipdriverout n19__chipdriverout 369e-3
rk20 n19__chipdriverout n20__chipdriverout 226.6e-3
rk21 n20__chipdriverout n21__chipdriverout 114.8e-3
rk22 n21__chipdriverout n22__chipdriverout 367.4e-3
rk23 n22__chipdriverout n23__chipdriverout 242.8e-3
rk24 n23__chipdriverout n24__chipdriverout 121.3e-3
rk26 n16__chipdriverout n17__chipdriverout 5.7692
rk27 n16__chipdriverout n20__chipdriverout 3.75
rk28 n16__chipdriverout n23__chipdriverout 3.75
rk29 n2__i1__i14__net1 n61__i1__i14__net1 125e-3
rk30 n4__i1__i14__net1 n62__i1__i14__net1 125e-3
rk31 n2__vss n3__vss 55.24e-3
rk32 n3__vss n4__vss 365.7e-3
rk33 n4__vss n5__vss 298.6e-3
rk34 n5__vss n6__vss 42.68e-3
rk35 n6__vss n7__vss 365.7e-3
rk36 n7__vss n8__vss 187.7e-3
rk37 n8__vss n9__vss 264.6e-3
rk38 n1__vss n2__vss 3.75
rk39 n1__vss n5__vss 3.75
rk40 n1__vss n8__vss 5.7692
rk42 n2__vddio n4__vddio 30.13e-3
rk43 n4__vddio n5__vddio 335.6e-3
rk44 n5__vddio n6__vddio 343.1e-3
rk45 n6__vddio n7__vddio 42.68e-3
rk46 n7__vddio n8__vddio 321.2e-3
rk47 n8__vddio n9__vddio 362.5e-3
rk48 n9__vddio n10__vddio 40.17e-3
rk49 n10__vddio n11__vddio 323.7e-3
rk50 n11__vddio n12__vddio 343.1e-3
rk51 n12__vddio n13__vddio 52.73e-3
rk52 n13__vddio n14__vddio 394.2e-3
rk53 n3__vddio n4__vddio 3.1
rk54 n3__vddio n7__vddio 3.1
rk55 n3__vddio n10__vddio 3.1
rk56 n3__vddio n13__vddio 3.1
rk57 n6__i1__i14__net1 n69__i1__i14__net1 125e-3
rk58 n8__i1__i14__net1 n70__i1__i14__net1 125e-3
rk60 n40__chipdriverout n42__chipdriverout 210.4e-3
rk61 n42__chipdriverout n43__chipdriverout 155.3e-3
rk62 n43__chipdriverout n44__chipdriverout 343.1e-3
rk63 n44__chipdriverout n45__chipdriverout 226.6e-3
rk64 n45__chipdriverout n46__chipdriverout 139.1e-3
rk65 n46__chipdriverout n47__chipdriverout 362.5e-3
rk66 n47__chipdriverout n48__chipdriverout 223.4e-3
rk67 n48__chipdriverout n49__chipdriverout 142.4e-3
rk68 n49__chipdriverout n50__chipdriverout 343.1e-3
rk69 n50__chipdriverout n51__chipdriverout 239.6e-3
rk70 n51__chipdriverout n52__chipdriverout 126.2e-3
rk72 n41__chipdriverout n42__chipdriverout 3.1
rk73 n41__chipdriverout n45__chipdriverout 3.1
rk74 n41__chipdriverout n48__chipdriverout 3.1
rk75 n41__chipdriverout n51__chipdriverout 3.1
rk77 n56__chipdriverout n57__chipdriverout 12.55e-3
rk78 n57__chipdriverout n58__chipdriverout 365.7e-3
rk79 n58__chipdriverout n59__chipdriverout 226.6e-3
rk80 n59__chipdriverout n60__chipdriverout 116.5e-3
rk81 n60__chipdriverout n61__chipdriverout 365.7e-3
rk82 n61__chipdriverout n62__chipdriverout 242.8e-3
rk83 n62__chipdriverout n63__chipdriverout 119.7e-3
rk85 n55__chipdriverout n56__chipdriverout 5.7692
rk86 n55__chipdriverout n59__chipdriverout 3.75
rk87 n55__chipdriverout n62__chipdriverout 3.75
rk88 n10__i1__i14__net1 n73__i1__i14__net1 125e-3
rk89 n12__i1__i14__net1 n74__i1__i14__net1 125e-3
rk90 n15__vss n16__vss 55.24e-3
rk91 n16__vss n17__vss 365.7e-3
rk92 n17__vss n18__vss 298.6e-3
rk93 n18__vss n19__vss 42.68e-3
rk94 n19__vss n20__vss 365.7e-3
rk95 n20__vss n21__vss 187.7e-3
rk96 n21__vss n22__vss 264.6e-3
rk97 n14__vss n15__vss 3.75
rk98 n14__vss n18__vss 3.75
rk99 n14__vss n21__vss 5.7692
rk101 n23__vddio n25__vddio 30.13e-3
rk102 n25__vddio n26__vddio 335.6e-3
rk103 n26__vddio n27__vddio 343.1e-3
rk104 n27__vddio n28__vddio 42.68e-3
rk105 n28__vddio n29__vddio 321.2e-3
rk106 n29__vddio n30__vddio 362.5e-3
rk107 n30__vddio n31__vddio 40.17e-3
rk108 n31__vddio n32__vddio 323.7e-3
rk109 n32__vddio n33__vddio 343.1e-3
rk110 n33__vddio n34__vddio 52.73e-3
rk111 n34__vddio n35__vddio 394.2e-3
rk112 n24__vddio n25__vddio 3.1
rk113 n24__vddio n28__vddio 3.1
rk114 n24__vddio n31__vddio 3.1
rk115 n24__vddio n34__vddio 3.1
rk119 n79__chipdriverout n81__chipdriverout 210.4e-3
rk120 n81__chipdriverout n82__chipdriverout 155.3e-3
rk121 n82__chipdriverout n83__chipdriverout 343.1e-3
rk122 n83__chipdriverout n84__chipdriverout 226.6e-3
rk123 n84__chipdriverout n85__chipdriverout 139.1e-3
rk124 n85__chipdriverout n86__chipdriverout 362.5e-3
rk125 n86__chipdriverout n87__chipdriverout 223.4e-3
rk126 n87__chipdriverout n88__chipdriverout 142.4e-3
rk127 n88__chipdriverout n89__chipdriverout 343.1e-3
rk128 n89__chipdriverout n90__chipdriverout 239.6e-3
rk129 n90__chipdriverout n91__chipdriverout 126.2e-3
rk131 n80__chipdriverout n81__chipdriverout 3.1
rk132 n80__chipdriverout n84__chipdriverout 3.1
rk133 n80__chipdriverout n87__chipdriverout 3.1
rk134 n80__chipdriverout n90__chipdriverout 3.1
rk136 n95__chipdriverout n96__chipdriverout 12.55e-3
rk137 n96__chipdriverout n97__chipdriverout 365.7e-3
rk138 n97__chipdriverout n98__chipdriverout 226.6e-3
rk139 n98__chipdriverout n99__chipdriverout 116.5e-3
rk140 n99__chipdriverout n100__chipdriverout 365.7e-3
rk141 n100__chipdriverout n101__chipdriverout 242.8e-3
rk142 n101__chipdriverout n102__chipdriverout 119.7e-3
rk144 n94__chipdriverout n95__chipdriverout 5.7692
rk145 n94__chipdriverout n98__chipdriverout 3.75
rk146 n94__chipdriverout n101__chipdriverout 3.75
rk147 n18__i1__i14__net1 n93__i1__i14__net1 125e-3
rk148 n20__i1__i14__net1 n94__i1__i14__net1 125e-3
rk149 n28__vss n29__vss 55.24e-3
rk150 n29__vss n30__vss 365.7e-3
rk151 n30__vss n31__vss 298.6e-3
rk152 n31__vss n32__vss 42.68e-3
rk153 n32__vss n33__vss 365.7e-3
rk154 n33__vss n34__vss 187.7e-3
rk155 n34__vss n35__vss 264.6e-3
rk156 n27__vss n28__vss 3.75
rk157 n27__vss n31__vss 3.75
rk158 n27__vss n34__vss 5.7692
rk160 n44__vddio n46__vddio 30.13e-3
rk161 n46__vddio n47__vddio 335.6e-3
rk162 n47__vddio n48__vddio 343.1e-3
rk163 n48__vddio n49__vddio 42.68e-3
rk164 n49__vddio n50__vddio 321.2e-3
rk165 n50__vddio n51__vddio 362.5e-3
rk166 n51__vddio n52__vddio 40.17e-3
rk167 n52__vddio n53__vddio 323.7e-3
rk168 n53__vddio n54__vddio 343.1e-3
rk169 n54__vddio n55__vddio 52.73e-3
rk170 n55__vddio n56__vddio 394.2e-3
rk171 n45__vddio n46__vddio 3.1
rk172 n45__vddio n49__vddio 3.1
rk173 n45__vddio n52__vddio 3.1
rk174 n45__vddio n55__vddio 3.1
rk175 n2__i5__clk4 n22__i5__clk4 45.506
rk176 n5__i5__clk4 n23__i5__clk4 45.506
rk177 n21__i1__i14__net1 n101__i1__i14__net1 125e-3
rk178 n23__i1__i14__net1 n102__i1__i14__net1 125e-3
rk179 n7__i5__i7__i0__net1 n8__i5__i7__i0__net1 75.2173
rk180 n7__i5__i7__i0__net1 n9__i5__i7__i0__net1 31.1536
rk181 n7__i5__i7__i1__net1 n8__i5__i7__i1__net1 75.2173
rk182 n7__i5__i7__i1__net1 n9__i5__i7__i1__net1 31.1536
rk184 n118__chipdriverout n120__chipdriverout 210.4e-3
rk185 n120__chipdriverout n121__chipdriverout 155.3e-3
rk186 n121__chipdriverout n122__chipdriverout 343.1e-3
rk187 n122__chipdriverout n123__chipdriverout 226.6e-3
rk188 n123__chipdriverout n124__chipdriverout 139.1e-3
rk189 n124__chipdriverout n125__chipdriverout 362.5e-3
rk190 n125__chipdriverout n126__chipdriverout 223.4e-3
rk191 n126__chipdriverout n127__chipdriverout 142.4e-3
rk192 n127__chipdriverout n128__chipdriverout 343.1e-3
rk193 n128__chipdriverout n129__chipdriverout 239.6e-3
rk194 n129__chipdriverout n130__chipdriverout 126.2e-3
rk196 n119__chipdriverout n120__chipdriverout 3.1
rk197 n119__chipdriverout n123__chipdriverout 3.1
rk198 n119__chipdriverout n126__chipdriverout 3.1
rk199 n119__chipdriverout n129__chipdriverout 3.1
rk201 n134__chipdriverout n135__chipdriverout 12.55e-3
rk202 n135__chipdriverout n136__chipdriverout 365.7e-3
rk203 n136__chipdriverout n137__chipdriverout 226.6e-3
rk204 n137__chipdriverout n138__chipdriverout 116.5e-3
rk205 n138__chipdriverout n139__chipdriverout 365.7e-3
rk206 n139__chipdriverout n140__chipdriverout 242.8e-3
rk207 n140__chipdriverout n141__chipdriverout 119.7e-3
rk209 n133__chipdriverout n134__chipdriverout 5.7692
rk210 n133__chipdriverout n137__chipdriverout 3.75
rk211 n133__chipdriverout n140__chipdriverout 3.75
rk212 n26__i1__i14__net1 n109__i1__i14__net1 125e-3
rk213 n28__i1__i14__net1 n110__i1__i14__net1 125e-3
rk214 n41__vss n42__vss 55.24e-3
rk215 n42__vss n43__vss 365.7e-3
rk216 n43__vss n44__vss 298.6e-3
rk217 n44__vss n45__vss 42.68e-3
rk218 n45__vss n46__vss 365.7e-3
rk219 n46__vss n47__vss 187.7e-3
rk220 n47__vss n48__vss 264.6e-3
rk221 n40__vss n41__vss 3.75
rk222 n40__vss n44__vss 3.75
rk223 n40__vss n47__vss 5.7692
rk225 n69__vddio n71__vddio 30.13e-3
rk226 n71__vddio n72__vddio 335.6e-3
rk227 n72__vddio n73__vddio 343.1e-3
rk228 n73__vddio n74__vddio 42.68e-3
rk229 n74__vddio n75__vddio 321.2e-3
rk230 n75__vddio n76__vddio 362.5e-3
rk231 n76__vddio n77__vddio 40.17e-3
rk232 n77__vddio n78__vddio 323.7e-3
rk233 n78__vddio n79__vddio 343.1e-3
rk234 n79__vddio n80__vddio 52.73e-3
rk235 n80__vddio n81__vddio 394.2e-3
rk236 n70__vddio n71__vddio 3.1
rk237 n70__vddio n74__vddio 3.1
rk238 n70__vddio n77__vddio 3.1
rk239 n70__vddio n80__vddio 3.1
rk241 n6__x0 n3__x0 4.923e-3
rk243 n6__y0 n3__y0 4.923e-3
rk244 n29__i1__i14__net1 n117__i1__i14__net1 125e-3
rk245 n31__i1__i14__net1 n118__i1__i14__net1 125e-3
rk247 n158__chipdriverout n159__chipdriverout 12.55e-3
rk248 n159__chipdriverout n160__chipdriverout 365.7e-3
rk249 n160__chipdriverout n161__chipdriverout 226.6e-3
rk250 n161__chipdriverout n162__chipdriverout 116.5e-3
rk251 n162__chipdriverout n163__chipdriverout 365.7e-3
rk252 n163__chipdriverout n164__chipdriverout 242.8e-3
rk253 n164__chipdriverout n165__chipdriverout 119.7e-3
rk255 n157__chipdriverout n158__chipdriverout 5.7692
rk256 n157__chipdriverout n161__chipdriverout 3.75
rk257 n157__chipdriverout n164__chipdriverout 3.75
rk259 n168__chipdriverout n170__chipdriverout 210.4e-3
rk260 n170__chipdriverout n171__chipdriverout 155.3e-3
rk261 n171__chipdriverout n172__chipdriverout 343.1e-3
rk262 n172__chipdriverout n173__chipdriverout 226.6e-3
rk263 n173__chipdriverout n174__chipdriverout 139.1e-3
rk264 n174__chipdriverout n175__chipdriverout 362.5e-3
rk265 n175__chipdriverout n176__chipdriverout 223.4e-3
rk266 n176__chipdriverout n177__chipdriverout 142.4e-3
rk267 n177__chipdriverout n178__chipdriverout 343.1e-3
rk268 n178__chipdriverout n179__chipdriverout 239.6e-3
rk269 n179__chipdriverout n180__chipdriverout 126.2e-3
rk271 n169__chipdriverout n170__chipdriverout 3.1
rk272 n169__chipdriverout n173__chipdriverout 3.1
rk273 n169__chipdriverout n176__chipdriverout 3.1
rk274 n169__chipdriverout n179__chipdriverout 3.1
rk277 i5__i7__i0__i3__net21 n2__i5__i7__i0__i3__net21 62.1844
rk278 i5__i7__i0__i3__net23 n2__i5__i7__i0__i3__net23 150.195
rk279 i5__i7__i1__i3__net21 n2__i5__i7__i1__i3__net21 62.1844
rk280 i5__i7__i1__i3__net23 n2__i5__i7__i1__i3__net23 150.195
rk281 n30__i5__clk4 n8__i5__clk4 505.3e-3
rk282 n13__i5__i7__i0__net1 n2__i5__i7__i0__net1 505.3e-3
rk283 n31__i5__clk4 n10__i5__clk4 505.3e-3
rk284 n13__i5__i7__i1__net1 n2__i5__i7__i1__net1 505.3e-3
rk285 n54__vss n55__vss 55.24e-3
rk286 n55__vss n56__vss 365.7e-3
rk287 n56__vss n57__vss 298.6e-3
rk288 n57__vss n58__vss 42.68e-3
rk289 n58__vss n59__vss 365.7e-3
rk290 n59__vss n60__vss 187.7e-3
rk291 n60__vss n61__vss 264.6e-3
rk292 n53__vss n54__vss 3.75
rk293 n53__vss n57__vss 3.75
rk294 n53__vss n60__vss 5.7692
rk296 n96__vddio n98__vddio 30.13e-3
rk297 n98__vddio n99__vddio 335.6e-3
rk298 n99__vddio n100__vddio 343.1e-3
rk299 n100__vddio n101__vddio 42.68e-3
rk300 n101__vddio n102__vddio 321.2e-3
rk301 n102__vddio n103__vddio 362.5e-3
rk302 n103__vddio n104__vddio 40.17e-3
rk303 n104__vddio n105__vddio 323.7e-3
rk304 n105__vddio n106__vddio 343.1e-3
rk305 n106__vddio n107__vddio 52.73e-3
rk306 n107__vddio n108__vddio 394.2e-3
rk307 n97__vddio n98__vddio 3.1
rk308 n97__vddio n101__vddio 3.1
rk309 n97__vddio n104__vddio 3.1
rk310 n97__vddio n107__vddio 3.1
rk311 n37__i1__i14__net1 n129__i1__i14__net1 125e-3
rk312 n39__i1__i14__net1 n130__i1__i14__net1 125e-3
rk314 n197__chipdriverout n198__chipdriverout 12.55e-3
rk315 n198__chipdriverout n199__chipdriverout 365.7e-3
rk316 n199__chipdriverout n200__chipdriverout 226.6e-3
rk317 n200__chipdriverout n201__chipdriverout 116.5e-3
rk318 n201__chipdriverout n202__chipdriverout 365.7e-3
rk319 n202__chipdriverout n203__chipdriverout 242.8e-3
rk320 n203__chipdriverout n204__chipdriverout 119.7e-3
rk322 n196__chipdriverout n197__chipdriverout 5.7692
rk323 n196__chipdriverout n200__chipdriverout 3.75
rk324 n196__chipdriverout n203__chipdriverout 3.75
rk326 n207__chipdriverout n209__chipdriverout 210.4e-3
rk327 n209__chipdriverout n210__chipdriverout 155.3e-3
rk328 n210__chipdriverout n211__chipdriverout 343.1e-3
rk329 n211__chipdriverout n212__chipdriverout 226.6e-3
rk330 n212__chipdriverout n213__chipdriverout 139.1e-3
rk331 n213__chipdriverout n214__chipdriverout 362.5e-3
rk332 n214__chipdriverout n215__chipdriverout 223.4e-3
rk333 n215__chipdriverout n216__chipdriverout 142.4e-3
rk334 n216__chipdriverout n217__chipdriverout 343.1e-3
rk335 n217__chipdriverout n218__chipdriverout 239.6e-3
rk336 n218__chipdriverout n219__chipdriverout 126.2e-3
rk338 n208__chipdriverout n209__chipdriverout 3.1
rk339 n208__chipdriverout n212__chipdriverout 3.1
rk340 n208__chipdriverout n215__chipdriverout 3.1
rk341 n208__chipdriverout n218__chipdriverout 3.1
rk342 n42__i1__i14__net1 n137__i1__i14__net1 125e-3
rk343 n44__i1__i14__net1 n138__i1__i14__net1 125e-3
rk344 n5__i5__i7__i0__i3__net22 n6__i5__i7__i0__i3__net22 31.2679
rk345 n6__i5__i7__i0__i3__net22 n7__i5__i7__i0__i3__net22 75.2632
rk346 n6__i5__i7__i0__i3__net22 n3__i5__i7__i0__i3__net22 230.1e-3
rk347 n5__i5__i7__i1__i3__net22 n6__i5__i7__i1__i3__net22 31.2679
rk348 n6__i5__i7__i1__i3__net22 n7__i5__i7__i1__i3__net22 75.2632
rk349 n6__i5__i7__i1__i3__net22 n3__i5__i7__i1__i3__net22 230.1e-3
rk351 n117__vddio n119__vddio 30.13e-3
rk352 n119__vddio n120__vddio 335.6e-3
rk353 n120__vddio n121__vddio 343.1e-3
rk354 n121__vddio n122__vddio 42.68e-3
rk355 n122__vddio n123__vddio 321.2e-3
rk356 n123__vddio n124__vddio 362.5e-3
rk357 n124__vddio n125__vddio 40.17e-3
rk358 n125__vddio n126__vddio 323.7e-3
rk359 n126__vddio n127__vddio 343.1e-3
rk360 n127__vddio n128__vddio 52.73e-3
rk361 n128__vddio n129__vddio 394.2e-3
rk362 n118__vddio n119__vddio 3.1
rk363 n118__vddio n122__vddio 3.1
rk364 n118__vddio n125__vddio 3.1
rk365 n118__vddio n128__vddio 3.1
rk366 n67__vss n68__vss 55.24e-3
rk367 n68__vss n69__vss 365.7e-3
rk368 n69__vss n70__vss 298.6e-3
rk369 n70__vss n71__vss 42.68e-3
rk370 n71__vss n72__vss 365.7e-3
rk371 n72__vss n73__vss 187.7e-3
rk372 n73__vss n74__vss 264.6e-3
rk373 n66__vss n67__vss 3.75
rk374 n66__vss n70__vss 3.75
rk375 n66__vss n73__vss 5.7692
rk376 n45__i1__i14__net1 n149__i1__i14__net1 125e-3
rk377 n47__i1__i14__net1 n150__i1__i14__net1 125e-3
rk378 i5__i7__i0__i3__net24 n2__i5__i7__i0__i3__net24 62.1844
rk379 i5__i7__i0__i3__net25 n2__i5__i7__i0__i3__net25 150.195
rk381 n236__chipdriverout n237__chipdriverout 12.55e-3
rk382 n237__chipdriverout n238__chipdriverout 365.7e-3
rk383 n238__chipdriverout n239__chipdriverout 226.6e-3
rk384 n239__chipdriverout n240__chipdriverout 116.5e-3
rk385 n240__chipdriverout n241__chipdriverout 365.7e-3
rk386 n241__chipdriverout n242__chipdriverout 242.8e-3
rk387 n242__chipdriverout n243__chipdriverout 119.7e-3
rk389 n235__chipdriverout n236__chipdriverout 5.7692
rk390 n235__chipdriverout n239__chipdriverout 3.75
rk391 n235__chipdriverout n242__chipdriverout 3.75
rk393 n246__chipdriverout n248__chipdriverout 210.4e-3
rk394 n248__chipdriverout n249__chipdriverout 155.3e-3
rk395 n249__chipdriverout n250__chipdriverout 343.1e-3
rk396 n250__chipdriverout n251__chipdriverout 226.6e-3
rk397 n251__chipdriverout n252__chipdriverout 139.1e-3
rk398 n252__chipdriverout n253__chipdriverout 362.5e-3
rk399 n253__chipdriverout n254__chipdriverout 223.4e-3
rk400 n254__chipdriverout n255__chipdriverout 142.4e-3
rk401 n255__chipdriverout n256__chipdriverout 343.1e-3
rk402 n256__chipdriverout n257__chipdriverout 239.6e-3
rk403 n257__chipdriverout n258__chipdriverout 126.2e-3
rk405 n247__chipdriverout n248__chipdriverout 3.1
rk406 n247__chipdriverout n251__chipdriverout 3.1
rk407 n247__chipdriverout n254__chipdriverout 3.1
rk408 n247__chipdriverout n257__chipdriverout 3.1
rk409 i5__i7__i1__i3__net24 n2__i5__i7__i1__i3__net24 62.1844
rk410 i5__i7__i1__i3__net25 n2__i5__i7__i1__i3__net25 150.195
rk411 n12__i5__clk4 n32__i5__clk4 4.923e-3
rk412 n14__i5__i7__i0__net1 n4__i5__i7__i0__net1 507.7e-3
rk413 n14__i5__clk4 n33__i5__clk4 4.923e-3
rk414 n14__i5__i7__i1__net1 n4__i5__i7__i1__net1 507.7e-3
rk415 n50__i1__i14__net1 n153__i1__i14__net1 125e-3
rk416 n52__i1__i14__net1 n154__i1__i14__net1 125e-3
rk418 n138__vddio n140__vddio 30.13e-3
rk419 n140__vddio n141__vddio 335.6e-3
rk420 n141__vddio n142__vddio 343.1e-3
rk421 n142__vddio n143__vddio 42.68e-3
rk422 n143__vddio n144__vddio 321.2e-3
rk423 n144__vddio n145__vddio 362.5e-3
rk424 n145__vddio n146__vddio 40.17e-3
rk425 n146__vddio n147__vddio 323.7e-3
rk426 n147__vddio n148__vddio 343.1e-3
rk427 n148__vddio n149__vddio 52.73e-3
rk428 n149__vddio n150__vddio 394.2e-3
rk429 n139__vddio n140__vddio 3.1
rk430 n139__vddio n143__vddio 3.1
rk431 n139__vddio n146__vddio 3.1
rk432 n139__vddio n149__vddio 3.1
rk433 n80__vss n81__vss 55.24e-3
rk434 n81__vss n82__vss 365.7e-3
rk435 n82__vss n83__vss 298.6e-3
rk436 n83__vss n84__vss 42.68e-3
rk437 n84__vss n85__vss 365.7e-3
rk438 n85__vss n86__vss 187.7e-3
rk439 n86__vss n87__vss 264.6e-3
rk440 n79__vss n80__vss 3.75
rk441 n79__vss n83__vss 3.75
rk442 n79__vss n86__vss 5.7692
rk443 n53__i1__i14__net1 n165__i1__i14__net1 125e-3
rk444 n55__i1__i14__net1 n166__i1__i14__net1 125e-3
rk445 n2__reset n9__reset 577.1e-3
rk446 n4__reset n12__reset 77.13e-3
rk448 n275__chipdriverout n276__chipdriverout 12.55e-3
rk449 n276__chipdriverout n277__chipdriverout 365.7e-3
rk450 n277__chipdriverout n278__chipdriverout 226.6e-3
rk451 n278__chipdriverout n279__chipdriverout 116.5e-3
rk452 n279__chipdriverout n280__chipdriverout 365.7e-3
rk453 n280__chipdriverout n281__chipdriverout 242.8e-3
rk454 n281__chipdriverout n282__chipdriverout 119.7e-3
rk456 n274__chipdriverout n275__chipdriverout 5.7692
rk457 n274__chipdriverout n278__chipdriverout 3.75
rk458 n274__chipdriverout n281__chipdriverout 3.75
rk460 n285__chipdriverout n287__chipdriverout 210.4e-3
rk461 n287__chipdriverout n288__chipdriverout 155.3e-3
rk462 n288__chipdriverout n289__chipdriverout 343.1e-3
rk463 n289__chipdriverout n290__chipdriverout 226.6e-3
rk464 n290__chipdriverout n291__chipdriverout 139.1e-3
rk465 n291__chipdriverout n292__chipdriverout 362.5e-3
rk466 n292__chipdriverout n293__chipdriverout 223.4e-3
rk467 n293__chipdriverout n294__chipdriverout 142.4e-3
rk468 n294__chipdriverout n295__chipdriverout 343.1e-3
rk469 n295__chipdriverout n296__chipdriverout 239.6e-3
rk470 n296__chipdriverout n297__chipdriverout 126.2e-3
rk472 n286__chipdriverout n287__chipdriverout 3.1
rk473 n286__chipdriverout n290__chipdriverout 3.1
rk474 n286__chipdriverout n293__chipdriverout 3.1
rk475 n286__chipdriverout n296__chipdriverout 3.1
rk476 i5__i7__x0out n2__i5__i7__x0out 19.2986
rk477 n2__i5__i7__x0out n4__i5__i7__x0out 528.7e-3
rk478 n4__i5__i7__x0out n5__i5__i7__x0out 75.4978
rk479 n3__i5__i7__x0out n4__i5__i7__x0out 31
rk480 i5__i7__y0out n2__i5__i7__y0out 19.2986
rk481 n2__i5__i7__y0out n4__i5__i7__y0out 528.7e-3
rk482 n4__i5__i7__y0out n5__i5__i7__y0out 75.4978
rk483 n3__i5__i7__y0out n4__i5__i7__y0out 31
rk487 n159__vddio n161__vddio 30.13e-3
rk488 n161__vddio n162__vddio 335.6e-3
rk489 n162__vddio n163__vddio 343.1e-3
rk490 n163__vddio n164__vddio 42.68e-3
rk491 n164__vddio n165__vddio 321.2e-3
rk492 n165__vddio n166__vddio 362.5e-3
rk493 n166__vddio n167__vddio 40.17e-3
rk494 n167__vddio n168__vddio 323.7e-3
rk495 n168__vddio n169__vddio 343.1e-3
rk496 n169__vddio n170__vddio 52.73e-3
rk497 n170__vddio n171__vddio 394.2e-3
rk498 n160__vddio n161__vddio 3.1
rk499 n160__vddio n164__vddio 3.1
rk500 n160__vddio n167__vddio 3.1
rk501 n160__vddio n170__vddio 3.1
rk502 n93__vss n94__vss 55.24e-3
rk503 n94__vss n95__vss 365.7e-3
rk504 n95__vss n96__vss 298.6e-3
rk505 n96__vss n97__vss 42.68e-3
rk506 n97__vss n98__vss 365.7e-3
rk507 n98__vss n99__vss 187.7e-3
rk508 n99__vss n100__vss 264.6e-3
rk509 n92__vss n93__vss 3.75
rk510 n92__vss n96__vss 3.75
rk511 n92__vss n99__vss 5.7692
rk512 n65__i1__i14__net1 n181__i1__i14__net1 125e-3
rk513 n67__i1__i14__net1 n182__i1__i14__net1 125e-3
rk515 n6__x1 n3__x1 4.923e-3
rk517 n7__y1 n3__y1 4.923e-3
rk519 n314__chipdriverout n315__chipdriverout 12.55e-3
rk520 n315__chipdriverout n316__chipdriverout 365.7e-3
rk521 n316__chipdriverout n317__chipdriverout 226.6e-3
rk522 n317__chipdriverout n318__chipdriverout 116.5e-3
rk523 n318__chipdriverout n319__chipdriverout 365.7e-3
rk524 n319__chipdriverout n320__chipdriverout 242.8e-3
rk525 n320__chipdriverout n321__chipdriverout 119.7e-3
rk527 n313__chipdriverout n314__chipdriverout 5.7692
rk528 n313__chipdriverout n317__chipdriverout 3.75
rk529 n313__chipdriverout n320__chipdriverout 3.75
rk531 n324__chipdriverout n326__chipdriverout 210.4e-3
rk532 n326__chipdriverout n327__chipdriverout 155.3e-3
rk533 n327__chipdriverout n328__chipdriverout 343.1e-3
rk534 n328__chipdriverout n329__chipdriverout 226.6e-3
rk535 n329__chipdriverout n330__chipdriverout 139.1e-3
rk536 n330__chipdriverout n331__chipdriverout 362.5e-3
rk537 n331__chipdriverout n332__chipdriverout 223.4e-3
rk538 n332__chipdriverout n333__chipdriverout 142.4e-3
rk539 n333__chipdriverout n334__chipdriverout 343.1e-3
rk540 n334__chipdriverout n335__chipdriverout 239.6e-3
rk541 n335__chipdriverout n336__chipdriverout 126.2e-3
rk543 n325__chipdriverout n326__chipdriverout 3.1
rk544 n325__chipdriverout n329__chipdriverout 3.1
rk545 n325__chipdriverout n332__chipdriverout 3.1
rk546 n325__chipdriverout n335__chipdriverout 3.1
rk547 n78__i1__i14__net1 n189__i1__i14__net1 125e-3
rk548 n80__i1__i14__net1 n190__i1__i14__net1 125e-3
rk550 n180__vddio n182__vddio 30.13e-3
rk551 n182__vddio n183__vddio 335.6e-3
rk552 n183__vddio n184__vddio 343.1e-3
rk553 n184__vddio n185__vddio 42.68e-3
rk554 n185__vddio n186__vddio 321.2e-3
rk555 n186__vddio n187__vddio 362.5e-3
rk556 n187__vddio n188__vddio 40.17e-3
rk557 n188__vddio n189__vddio 323.7e-3
rk558 n189__vddio n190__vddio 343.1e-3
rk559 n190__vddio n191__vddio 52.73e-3
rk560 n191__vddio n192__vddio 394.2e-3
rk561 n181__vddio n182__vddio 3.1
rk562 n181__vddio n185__vddio 3.1
rk563 n181__vddio n188__vddio 3.1
rk564 n181__vddio n191__vddio 3.1
rk565 n106__vss n107__vss 55.24e-3
rk566 n107__vss n108__vss 365.7e-3
rk567 n108__vss n109__vss 298.6e-3
rk568 n109__vss n110__vss 42.68e-3
rk569 n110__vss n111__vss 365.7e-3
rk570 n111__vss n112__vss 187.7e-3
rk571 n112__vss n113__vss 264.6e-3
rk572 n105__vss n106__vss 3.75
rk573 n105__vss n109__vss 3.75
rk574 n105__vss n112__vss 5.7692
rk575 i5__i7__i0__i0__net21 n2__i5__i7__i0__i0__net21 62.1844
rk576 i5__i7__i0__i0__net23 n2__i5__i7__i0__i0__net23 150.195
rk577 i5__i7__i1__i0__net21 n2__i5__i7__i1__i0__net21 62.1844
rk578 i5__i7__i1__i0__net23 n2__i5__i7__i1__i0__net23 150.195
rk579 n44__i5__clk4 n16__i5__clk4 505.3e-3
rk580 n20__i5__i7__i0__net1 n6__i5__i7__i0__net1 505.3e-3
rk583 n45__i5__clk4 n18__i5__clk4 505.3e-3
rk584 n20__i5__i7__i1__net1 n6__i5__i7__i1__net1 505.3e-3
rk586 n353__chipdriverout n354__chipdriverout 12.55e-3
rk587 n354__chipdriverout n355__chipdriverout 365.7e-3
rk588 n355__chipdriverout n356__chipdriverout 226.6e-3
rk589 n356__chipdriverout n357__chipdriverout 116.5e-3
rk590 n357__chipdriverout n358__chipdriverout 365.7e-3
rk591 n358__chipdriverout n359__chipdriverout 242.8e-3
rk592 n359__chipdriverout n360__chipdriverout 119.7e-3
rk594 n352__chipdriverout n353__chipdriverout 5.7692
rk595 n352__chipdriverout n356__chipdriverout 3.75
rk596 n352__chipdriverout n359__chipdriverout 3.75
rk598 n363__chipdriverout n365__chipdriverout 210.4e-3
rk599 n365__chipdriverout n366__chipdriverout 155.3e-3
rk600 n366__chipdriverout n367__chipdriverout 343.1e-3
rk601 n367__chipdriverout n368__chipdriverout 226.6e-3
rk602 n368__chipdriverout n369__chipdriverout 139.1e-3
rk603 n369__chipdriverout n370__chipdriverout 362.5e-3
rk604 n370__chipdriverout n371__chipdriverout 223.4e-3
rk605 n371__chipdriverout n372__chipdriverout 142.4e-3
rk606 n372__chipdriverout n373__chipdriverout 343.1e-3
rk607 n373__chipdriverout n374__chipdriverout 239.6e-3
rk608 n374__chipdriverout n375__chipdriverout 126.2e-3
rk610 n364__chipdriverout n365__chipdriverout 3.1
rk611 n364__chipdriverout n368__chipdriverout 3.1
rk612 n364__chipdriverout n371__chipdriverout 3.1
rk613 n364__chipdriverout n374__chipdriverout 3.1
rk617 n211__vddio n213__vddio 30.13e-3
rk618 n213__vddio n214__vddio 335.6e-3
rk619 n214__vddio n215__vddio 343.1e-3
rk620 n215__vddio n216__vddio 42.68e-3
rk621 n216__vddio n217__vddio 321.2e-3
rk622 n217__vddio n218__vddio 362.5e-3
rk623 n218__vddio n219__vddio 40.17e-3
rk624 n219__vddio n220__vddio 323.7e-3
rk625 n220__vddio n221__vddio 343.1e-3
rk626 n221__vddio n222__vddio 52.73e-3
rk627 n222__vddio n223__vddio 394.2e-3
rk628 n212__vddio n213__vddio 3.1
rk629 n212__vddio n216__vddio 3.1
rk630 n212__vddio n219__vddio 3.1
rk631 n212__vddio n222__vddio 3.1
rk632 n119__vss n120__vss 55.24e-3
rk633 n120__vss n121__vss 365.7e-3
rk634 n121__vss n122__vss 298.6e-3
rk635 n122__vss n123__vss 42.68e-3
rk636 n123__vss n124__vss 365.7e-3
rk637 n124__vss n125__vss 187.7e-3
rk638 n125__vss n126__vss 264.6e-3
rk639 n118__vss n119__vss 3.75
rk640 n118__vss n122__vss 3.75
rk641 n118__vss n125__vss 5.7692
rk642 n5__i5__i7__i0__i0__net22 n6__i5__i7__i0__i0__net22 31.2679
rk643 n6__i5__i7__i0__i0__net22 n7__i5__i7__i0__i0__net22 75.2632
rk644 n6__i5__i7__i0__i0__net22 n3__i5__i7__i0__i0__net22 230.1e-3
rk645 n5__i5__i7__i1__i0__net22 n6__i5__i7__i1__i0__net22 31.2679
rk646 n6__i5__i7__i1__i0__net22 n7__i5__i7__i1__i0__net22 75.2632
rk647 n6__i5__i7__i1__i0__net22 n3__i5__i7__i1__i0__net22 230.1e-3
rk648 n98__i1__i14__net1 n213__i1__i14__net1 125e-3
rk649 n100__i1__i14__net1 n214__i1__i14__net1 125e-3
rk651 n392__chipdriverout n393__chipdriverout 12.55e-3
rk652 n393__chipdriverout n394__chipdriverout 365.7e-3
rk653 n394__chipdriverout n395__chipdriverout 226.6e-3
rk654 n395__chipdriverout n396__chipdriverout 116.5e-3
rk655 n396__chipdriverout n397__chipdriverout 365.7e-3
rk656 n397__chipdriverout n398__chipdriverout 242.8e-3
rk657 n398__chipdriverout n399__chipdriverout 119.7e-3
rk659 n391__chipdriverout n392__chipdriverout 5.7692
rk660 n391__chipdriverout n395__chipdriverout 3.75
rk661 n391__chipdriverout n398__chipdriverout 3.75
rk663 n402__chipdriverout n404__chipdriverout 210.4e-3
rk664 n404__chipdriverout n405__chipdriverout 155.3e-3
rk665 n405__chipdriverout n406__chipdriverout 343.1e-3
rk666 n406__chipdriverout n407__chipdriverout 226.6e-3
rk667 n407__chipdriverout n408__chipdriverout 139.1e-3
rk668 n408__chipdriverout n409__chipdriverout 362.5e-3
rk669 n409__chipdriverout n410__chipdriverout 223.4e-3
rk670 n410__chipdriverout n411__chipdriverout 142.4e-3
rk671 n411__chipdriverout n412__chipdriverout 343.1e-3
rk672 n412__chipdriverout n413__chipdriverout 239.6e-3
rk673 n413__chipdriverout n414__chipdriverout 126.2e-3
rk675 n403__chipdriverout n404__chipdriverout 3.1
rk676 n403__chipdriverout n407__chipdriverout 3.1
rk677 n403__chipdriverout n410__chipdriverout 3.1
rk678 n403__chipdriverout n413__chipdriverout 3.1
rk679 n106__i1__i14__net1 n221__i1__i14__net1 125e-3
rk680 n108__i1__i14__net1 n222__i1__i14__net1 125e-3
rk681 i5__i7__i0__i0__net24 n2__i5__i7__i0__i0__net24 62.1844
rk682 i5__i7__i0__i0__net25 n2__i5__i7__i0__i0__net25 150.195
rk683 i5__i7__i1__i0__net24 n2__i5__i7__i1__i0__net24 62.1844
rk684 i5__i7__i1__i0__net25 n2__i5__i7__i1__i0__net25 150.195
rk685 n27__i5__clk4 n50__i5__clk4 4.923e-3
rk686 n23__i5__i7__i0__net1 n12__i5__i7__i0__net1 7.702e-3
rk687 n29__i5__clk4 n52__i5__clk4 4.923e-3
rk688 n23__i5__i7__i1__net1 n12__i5__i7__i1__net1 7.702e-3
rk690 n232__vddio n247__vddio 30.13e-3
rk691 n247__vddio n233__vddio 335.6e-3
rk692 n233__vddio n236__vddio 343.1e-3
rk693 n236__vddio n248__vddio 42.68e-3
rk694 n248__vddio n237__vddio 321.2e-3
rk695 n237__vddio n240__vddio 362.5e-3
rk696 n240__vddio n249__vddio 40.17e-3
rk697 n249__vddio n241__vddio 323.7e-3
rk698 n241__vddio n244__vddio 343.1e-3
rk699 n244__vddio n250__vddio 52.73e-3
rk700 n250__vddio n251__vddio 394.2e-3
rk701 n246__vddio n247__vddio 3.1
rk702 n246__vddio n248__vddio 3.1
rk703 n246__vddio n249__vddio 3.1
rk704 n246__vddio n250__vddio 3.1
rk705 n140__vss n137__vss 55.24e-3
rk706 n137__vss n136__vss 365.7e-3
rk707 n136__vss n141__vss 298.6e-3
rk708 n141__vss n133__vss 42.68e-3
rk709 n133__vss n132__vss 365.7e-3
rk710 n132__vss n142__vss 187.7e-3
rk711 n142__vss n143__vss 264.6e-3
rk712 n139__vss n140__vss 3.75
rk713 n139__vss n141__vss 3.75
rk714 n139__vss n142__vss 5.7692
rk715 n114__i1__i14__net1 n229__i1__i14__net1 125e-3
rk716 n116__i1__i14__net1 n230__i1__i14__net1 125e-3
rk718 n431__chipdriverout n432__chipdriverout 12.55e-3
rk719 n432__chipdriverout n433__chipdriverout 365.7e-3
rk720 n433__chipdriverout n434__chipdriverout 226.6e-3
rk721 n434__chipdriverout n435__chipdriverout 116.5e-3
rk722 n435__chipdriverout n436__chipdriverout 365.7e-3
rk723 n436__chipdriverout n437__chipdriverout 242.8e-3
rk724 n437__chipdriverout n438__chipdriverout 119.7e-3
rk726 n430__chipdriverout n431__chipdriverout 5.7692
rk727 n430__chipdriverout n434__chipdriverout 3.75
rk728 n430__chipdriverout n437__chipdriverout 3.75
rk730 n441__chipdriverout n443__chipdriverout 210.4e-3
rk731 n443__chipdriverout n444__chipdriverout 155.3e-3
rk732 n444__chipdriverout n445__chipdriverout 343.1e-3
rk733 n445__chipdriverout n446__chipdriverout 226.6e-3
rk734 n446__chipdriverout n447__chipdriverout 139.1e-3
rk735 n447__chipdriverout n448__chipdriverout 362.5e-3
rk736 n448__chipdriverout n449__chipdriverout 223.4e-3
rk737 n449__chipdriverout n450__chipdriverout 142.4e-3
rk738 n450__chipdriverout n451__chipdriverout 343.1e-3
rk739 n451__chipdriverout n452__chipdriverout 239.6e-3
rk740 n452__chipdriverout n453__chipdriverout 126.2e-3
rk742 n442__chipdriverout n443__chipdriverout 3.1
rk743 n442__chipdriverout n446__chipdriverout 3.1
rk744 n442__chipdriverout n449__chipdriverout 3.1
rk745 n442__chipdriverout n452__chipdriverout 3.1
rk746 n126__i1__i14__net1 n233__i1__i14__net1 125e-3
rk747 n128__i1__i14__net1 n234__i1__i14__net1 125e-3
rk748 n6__reset n20__reset 577.1e-3
rk749 n8__reset n21__reset 577.1e-3
rk751 n253__vddio n255__vddio 30.13e-3
rk752 n255__vddio n256__vddio 335.6e-3
rk753 n256__vddio n257__vddio 343.1e-3
rk754 n257__vddio n258__vddio 42.68e-3
rk755 n258__vddio n259__vddio 321.2e-3
rk756 n259__vddio n260__vddio 362.5e-3
rk757 n260__vddio n261__vddio 40.17e-3
rk758 n261__vddio n262__vddio 323.7e-3
rk759 n262__vddio n263__vddio 343.1e-3
rk760 n263__vddio n264__vddio 52.73e-3
rk761 n264__vddio n265__vddio 394.2e-3
rk762 n254__vddio n255__vddio 3.1
rk763 n254__vddio n258__vddio 3.1
rk764 n254__vddio n261__vddio 3.1
rk765 n254__vddio n264__vddio 3.1
rk766 n145__vss n146__vss 55.24e-3
rk767 n146__vss n147__vss 365.7e-3
rk768 n147__vss n148__vss 298.6e-3
rk769 n148__vss n149__vss 42.68e-3
rk770 n149__vss n150__vss 365.7e-3
rk771 n150__vss n151__vss 187.7e-3
rk772 n151__vss n152__vss 264.6e-3
rk773 n144__vss n145__vss 3.75
rk774 n144__vss n148__vss 3.75
rk775 n144__vss n151__vss 5.7692
rk776 i5__i7__x1out n2__i5__i7__x1out 19.2986
rk777 n2__i5__i7__x1out n4__i5__i7__x1out 528.7e-3
rk778 n4__i5__i7__x1out n5__i5__i7__x1out 75.4978
rk779 n3__i5__i7__x1out n4__i5__i7__x1out 31
rk780 i5__i7__y1out n2__i5__i7__y1out 19.2986
rk781 n2__i5__i7__y1out n4__i5__i7__y1out 528.7e-3
rk782 n4__i5__i7__y1out n5__i5__i7__y1out 75.4978
rk783 n3__i5__i7__y1out n4__i5__i7__y1out 31
rk784 n132__i1__i14__net1 n245__i1__i14__net1 125e-3
rk785 n134__i1__i14__net1 n246__i1__i14__net1 125e-3
rk787 n469__chipdriverout n471__chipdriverout 210.4e-3
rk788 n471__chipdriverout n472__chipdriverout 155.3e-3
rk789 n472__chipdriverout n473__chipdriverout 343.1e-3
rk790 n473__chipdriverout n474__chipdriverout 226.6e-3
rk791 n474__chipdriverout n475__chipdriverout 139.1e-3
rk792 n475__chipdriverout n476__chipdriverout 362.5e-3
rk793 n476__chipdriverout n477__chipdriverout 223.4e-3
rk794 n477__chipdriverout n478__chipdriverout 142.4e-3
rk795 n478__chipdriverout n479__chipdriverout 343.1e-3
rk796 n479__chipdriverout n480__chipdriverout 239.6e-3
rk797 n480__chipdriverout n481__chipdriverout 126.2e-3
rk799 n470__chipdriverout n471__chipdriverout 3.1
rk800 n470__chipdriverout n474__chipdriverout 3.1
rk801 n470__chipdriverout n477__chipdriverout 3.1
rk802 n470__chipdriverout n480__chipdriverout 3.1
rk804 n485__chipdriverout n486__chipdriverout 12.55e-3
rk805 n486__chipdriverout n487__chipdriverout 365.7e-3
rk806 n487__chipdriverout n488__chipdriverout 226.6e-3
rk807 n488__chipdriverout n489__chipdriverout 116.5e-3
rk808 n489__chipdriverout n490__chipdriverout 365.7e-3
rk809 n490__chipdriverout n491__chipdriverout 242.8e-3
rk810 n491__chipdriverout n492__chipdriverout 119.7e-3
rk812 n484__chipdriverout n485__chipdriverout 5.7692
rk813 n484__chipdriverout n488__chipdriverout 3.75
rk814 n484__chipdriverout n491__chipdriverout 3.75
rk816 n6__x2 n3__x2 4.923e-3
rk818 n6__y2 n3__y2 4.923e-3
rk822 n284__vddio n286__vddio 30.13e-3
rk823 n286__vddio n287__vddio 335.6e-3
rk824 n287__vddio n288__vddio 343.1e-3
rk825 n288__vddio n289__vddio 42.68e-3
rk826 n289__vddio n290__vddio 321.2e-3
rk827 n290__vddio n291__vddio 362.5e-3
rk828 n291__vddio n292__vddio 40.17e-3
rk829 n292__vddio n293__vddio 323.7e-3
rk830 n293__vddio n294__vddio 343.1e-3
rk831 n294__vddio n295__vddio 52.73e-3
rk832 n295__vddio n296__vddio 394.2e-3
rk833 n285__vddio n286__vddio 3.1
rk834 n285__vddio n289__vddio 3.1
rk835 n285__vddio n292__vddio 3.1
rk836 n285__vddio n295__vddio 3.1
rk837 n158__vss n159__vss 55.24e-3
rk838 n159__vss n160__vss 365.7e-3
rk839 n160__vss n161__vss 298.6e-3
rk840 n161__vss n162__vss 42.68e-3
rk841 n162__vss n163__vss 365.7e-3
rk842 n163__vss n164__vss 187.7e-3
rk843 n164__vss n165__vss 264.6e-3
rk844 n157__vss n158__vss 3.75
rk845 n157__vss n161__vss 3.75
rk846 n157__vss n164__vss 5.7692
rk847 n146__i1__i14__net1 n261__i1__i14__net1 125e-3
rk848 n148__i1__i14__net1 n262__i1__i14__net1 125e-3
rk849 i5__i7__i0__i1__net21 n2__i5__i7__i0__i1__net21 62.1844
rk850 i5__i7__i0__i1__net23 n2__i5__i7__i0__i1__net23 150.195
rk851 i5__i7__i1__i1__net21 n2__i5__i7__i1__i1__net21 62.1844
rk852 i5__i7__i1__i1__net23 n2__i5__i7__i1__i1__net23 150.195
rk854 n518__chipdriverout n535__chipdriverout 210.4e-3
rk855 n535__chipdriverout n519__chipdriverout 155.3e-3
rk856 n519__chipdriverout n522__chipdriverout 343.1e-3
rk857 n522__chipdriverout n536__chipdriverout 226.6e-3
rk858 n536__chipdriverout n523__chipdriverout 139.1e-3
rk859 n523__chipdriverout n526__chipdriverout 362.5e-3
rk860 n526__chipdriverout n537__chipdriverout 223.4e-3
rk861 n537__chipdriverout n527__chipdriverout 142.4e-3
rk862 n527__chipdriverout n530__chipdriverout 343.1e-3
rk863 n530__chipdriverout n538__chipdriverout 239.6e-3
rk864 n538__chipdriverout n531__chipdriverout 126.2e-3
rk866 n534__chipdriverout n535__chipdriverout 3.1
rk867 n534__chipdriverout n536__chipdriverout 3.1
rk868 n534__chipdriverout n537__chipdriverout 3.1
rk869 n534__chipdriverout n538__chipdriverout 3.1
rk871 n542__chipdriverout n507__chipdriverout 12.55e-3
rk872 n507__chipdriverout n510__chipdriverout 365.7e-3
rk873 n510__chipdriverout n543__chipdriverout 226.6e-3
rk874 n543__chipdriverout n511__chipdriverout 116.5e-3
rk875 n511__chipdriverout n514__chipdriverout 365.7e-3
rk876 n514__chipdriverout n544__chipdriverout 242.8e-3
rk877 n544__chipdriverout n515__chipdriverout 119.7e-3
rk879 n541__chipdriverout n542__chipdriverout 5.7692
rk880 n541__chipdriverout n543__chipdriverout 3.75
rk881 n541__chipdriverout n544__chipdriverout 3.75
rk882 n58__i5__clk4 n37__i5__clk4 505.3e-3
rk883 n27__i5__i7__i0__net1 n17__i5__i7__i0__net1 505.3e-3
rk884 n59__i5__clk4 n39__i5__clk4 505.3e-3
rk885 n27__i5__i7__i1__net1 n17__i5__i7__i1__net1 505.3e-3
rk886 n158__i1__i14__net1 n265__i1__i14__net1 125e-3
rk887 n160__i1__i14__net1 n266__i1__i14__net1 125e-3
rk889 n305__vddio n320__vddio 30.13e-3
rk890 n320__vddio n306__vddio 335.6e-3
rk891 n306__vddio n309__vddio 343.1e-3
rk892 n309__vddio n321__vddio 42.68e-3
rk893 n321__vddio n310__vddio 321.2e-3
rk894 n310__vddio n313__vddio 362.5e-3
rk895 n313__vddio n322__vddio 40.17e-3
rk896 n322__vddio n314__vddio 323.7e-3
rk897 n314__vddio n317__vddio 343.1e-3
rk898 n317__vddio n323__vddio 52.73e-3
rk899 n323__vddio n324__vddio 394.2e-3
rk900 n319__vddio n320__vddio 3.1
rk901 n319__vddio n321__vddio 3.1
rk902 n319__vddio n322__vddio 3.1
rk903 n319__vddio n323__vddio 3.1
rk904 n179__vss n176__vss 55.24e-3
rk905 n176__vss n175__vss 365.7e-3
rk906 n175__vss n180__vss 298.6e-3
rk907 n180__vss n172__vss 42.68e-3
rk908 n172__vss n171__vss 365.7e-3
rk909 n171__vss n181__vss 187.7e-3
rk910 n181__vss n182__vss 264.6e-3
rk911 n178__vss n179__vss 3.75
rk912 n178__vss n180__vss 3.75
rk913 n178__vss n181__vss 5.7692
rk916 n5__i5__i7__i0__i1__net22 n6__i5__i7__i0__i1__net22 31.2679
rk917 n6__i5__i7__i0__i1__net22 n7__i5__i7__i0__i1__net22 75.2632
rk918 n6__i5__i7__i0__i1__net22 n3__i5__i7__i0__i1__net22 230.1e-3
rk919 n5__i5__i7__i1__i1__net22 n6__i5__i7__i1__i1__net22 31.2679
rk920 n6__i5__i7__i1__i1__net22 n7__i5__i7__i1__i1__net22 75.2632
rk921 n6__i5__i7__i1__i1__net22 n3__i5__i7__i1__i1__net22 230.1e-3
rk923 n557__chipdriverout n574__chipdriverout 210.4e-3
rk924 n574__chipdriverout n558__chipdriverout 155.3e-3
rk925 n558__chipdriverout n561__chipdriverout 343.1e-3
rk926 n561__chipdriverout n575__chipdriverout 226.6e-3
rk927 n575__chipdriverout n562__chipdriverout 139.1e-3
rk928 n562__chipdriverout n565__chipdriverout 362.5e-3
rk929 n565__chipdriverout n576__chipdriverout 223.4e-3
rk930 n576__chipdriverout n566__chipdriverout 142.4e-3
rk931 n566__chipdriverout n569__chipdriverout 343.1e-3
rk932 n569__chipdriverout n577__chipdriverout 239.6e-3
rk933 n577__chipdriverout n570__chipdriverout 126.2e-3
rk935 n573__chipdriverout n574__chipdriverout 3.1
rk936 n573__chipdriverout n575__chipdriverout 3.1
rk937 n573__chipdriverout n576__chipdriverout 3.1
rk938 n573__chipdriverout n577__chipdriverout 3.1
rk940 n581__chipdriverout n546__chipdriverout 12.55e-3
rk941 n546__chipdriverout n549__chipdriverout 365.7e-3
rk942 n549__chipdriverout n582__chipdriverout 226.6e-3
rk943 n582__chipdriverout n550__chipdriverout 116.5e-3
rk944 n550__chipdriverout n553__chipdriverout 365.7e-3
rk945 n553__chipdriverout n583__chipdriverout 242.8e-3
rk946 n583__chipdriverout n554__chipdriverout 119.7e-3
rk948 n580__chipdriverout n581__chipdriverout 5.7692
rk949 n580__chipdriverout n582__chipdriverout 3.75
rk950 n580__chipdriverout n583__chipdriverout 3.75
rk951 n174__i1__i14__net1 n281__i1__i14__net1 125e-3
rk952 n176__i1__i14__net1 n282__i1__i14__net1 125e-3
rk954 n326__vddio n328__vddio 30.13e-3
rk955 n328__vddio n329__vddio 335.6e-3
rk956 n329__vddio n330__vddio 343.1e-3
rk957 n330__vddio n331__vddio 42.68e-3
rk958 n331__vddio n332__vddio 321.2e-3
rk959 n332__vddio n333__vddio 362.5e-3
rk960 n333__vddio n334__vddio 40.17e-3
rk961 n334__vddio n335__vddio 323.7e-3
rk962 n335__vddio n336__vddio 343.1e-3
rk963 n336__vddio n337__vddio 52.73e-3
rk964 n337__vddio n338__vddio 394.2e-3
rk965 n327__vddio n328__vddio 3.1
rk966 n327__vddio n331__vddio 3.1
rk967 n327__vddio n334__vddio 3.1
rk968 n327__vddio n337__vddio 3.1
rk969 n184__vss n185__vss 55.24e-3
rk970 n185__vss n186__vss 365.7e-3
rk971 n186__vss n187__vss 298.6e-3
rk972 n187__vss n188__vss 42.68e-3
rk973 n188__vss n189__vss 365.7e-3
rk974 n189__vss n190__vss 187.7e-3
rk975 n190__vss n191__vss 264.6e-3
rk976 n183__vss n184__vss 3.75
rk977 n183__vss n187__vss 3.75
rk978 n183__vss n190__vss 5.7692
rk979 i5__i7__i0__i1__net24 n2__i5__i7__i0__i1__net24 62.1844
rk980 i5__i7__i0__i1__net25 n2__i5__i7__i0__i1__net25 150.195
rk981 i5__i7__i1__i1__net24 n2__i5__i7__i1__i1__net24 62.1844
rk982 i5__i7__i1__i1__net25 n2__i5__i7__i1__i1__net25 150.195
rk983 n41__i5__clk4 n60__i5__clk4 4.923e-3
rk984 n28__i5__i7__i0__net1 n19__i5__i7__i0__net1 507.7e-3
rk985 n43__i5__clk4 n61__i5__clk4 4.923e-3
rk986 n28__i5__i7__i1__net1 n19__i5__i7__i1__net1 507.7e-3
rk987 n178__i1__i14__net1 n289__i1__i14__net1 125e-3
rk988 n180__i1__i14__net1 n290__i1__i14__net1 125e-3
rk990 n586__chipdriverout n588__chipdriverout 210.4e-3
rk991 n588__chipdriverout n589__chipdriverout 155.3e-3
rk992 n589__chipdriverout n590__chipdriverout 343.1e-3
rk993 n590__chipdriverout n591__chipdriverout 226.6e-3
rk994 n591__chipdriverout n592__chipdriverout 139.1e-3
rk995 n592__chipdriverout n593__chipdriverout 362.5e-3
rk996 n593__chipdriverout n594__chipdriverout 223.4e-3
rk997 n594__chipdriverout n595__chipdriverout 142.4e-3
rk998 n595__chipdriverout n596__chipdriverout 343.1e-3
rk999 n596__chipdriverout n597__chipdriverout 239.6e-3
rk1000 n597__chipdriverout n598__chipdriverout 126.2e-3
rk1002 n587__chipdriverout n588__chipdriverout 3.1
rk1003 n587__chipdriverout n591__chipdriverout 3.1
rk1004 n587__chipdriverout n594__chipdriverout 3.1
rk1005 n587__chipdriverout n597__chipdriverout 3.1
rk1007 n602__chipdriverout n603__chipdriverout 12.55e-3
rk1008 n603__chipdriverout n604__chipdriverout 365.7e-3
rk1009 n604__chipdriverout n605__chipdriverout 226.6e-3
rk1010 n605__chipdriverout n606__chipdriverout 116.5e-3
rk1011 n606__chipdriverout n607__chipdriverout 365.7e-3
rk1012 n607__chipdriverout n608__chipdriverout 242.8e-3
rk1013 n608__chipdriverout n609__chipdriverout 119.7e-3
rk1015 n601__chipdriverout n602__chipdriverout 5.7692
rk1016 n601__chipdriverout n605__chipdriverout 3.75
rk1017 n601__chipdriverout n608__chipdriverout 3.75
rk1020 n17__reset n29__reset 77.13e-3
rk1022 n347__vddio n362__vddio 30.13e-3
rk1023 n362__vddio n348__vddio 335.6e-3
rk1024 n348__vddio n351__vddio 343.1e-3
rk1025 n351__vddio n363__vddio 42.68e-3
rk1026 n363__vddio n352__vddio 321.2e-3
rk1027 n352__vddio n355__vddio 362.5e-3
rk1028 n355__vddio n364__vddio 40.17e-3
rk1029 n364__vddio n356__vddio 323.7e-3
rk1030 n356__vddio n359__vddio 343.1e-3
rk1031 n359__vddio n365__vddio 52.73e-3
rk1032 n365__vddio n366__vddio 394.2e-3
rk1033 n361__vddio n362__vddio 3.1
rk1034 n361__vddio n363__vddio 3.1
rk1035 n361__vddio n364__vddio 3.1
rk1036 n361__vddio n365__vddio 3.1
rk1037 n205__vss n202__vss 55.24e-3
rk1038 n202__vss n201__vss 365.7e-3
rk1039 n201__vss n206__vss 298.6e-3
rk1040 n206__vss n198__vss 42.68e-3
rk1041 n198__vss n197__vss 365.7e-3
rk1042 n197__vss n207__vss 187.7e-3
rk1043 n207__vss n208__vss 264.6e-3
rk1044 n204__vss n205__vss 3.75
rk1045 n204__vss n206__vss 3.75
rk1046 n204__vss n207__vss 5.7692
rk1047 n19__reset n31__reset 77.13e-3
rk1048 n4__i5__i7__x2out n5__i5__i7__x2out 19.2986
rk1049 n5__i5__i7__x2out n7__i5__i7__x2out 528.7e-3
rk1050 n7__i5__i7__x2out n8__i5__i7__x2out 75.4978
rk1051 n6__i5__i7__x2out n7__i5__i7__x2out 31
rk1052 n4__i5__i7__y2out n5__i5__i7__y2out 19.2986
rk1053 n5__i5__i7__y2out n7__i5__i7__y2out 528.7e-3
rk1054 n7__i5__i7__y2out n8__i5__i7__y2out 75.4978
rk1055 n6__i5__i7__y2out n7__i5__i7__y2out 31
rk1056 n198__i1__i14__net1 n309__i1__i14__net1 125e-3
rk1057 n200__i1__i14__net1 n310__i1__i14__net1 125e-3
rk1059 n625__chipdriverout n627__chipdriverout 210.4e-3
rk1060 n627__chipdriverout n628__chipdriverout 155.3e-3
rk1061 n628__chipdriverout n629__chipdriverout 343.1e-3
rk1062 n629__chipdriverout n630__chipdriverout 226.6e-3
rk1063 n630__chipdriverout n631__chipdriverout 139.1e-3
rk1064 n631__chipdriverout n632__chipdriverout 362.5e-3
rk1065 n632__chipdriverout n633__chipdriverout 223.4e-3
rk1066 n633__chipdriverout n634__chipdriverout 142.4e-3
rk1067 n634__chipdriverout n635__chipdriverout 343.1e-3
rk1068 n635__chipdriverout n636__chipdriverout 239.6e-3
rk1069 n636__chipdriverout n637__chipdriverout 126.2e-3
rk1071 n626__chipdriverout n627__chipdriverout 3.1
rk1072 n626__chipdriverout n630__chipdriverout 3.1
rk1073 n626__chipdriverout n633__chipdriverout 3.1
rk1074 n626__chipdriverout n636__chipdriverout 3.1
rk1076 n641__chipdriverout n642__chipdriverout 12.55e-3
rk1077 n642__chipdriverout n643__chipdriverout 365.7e-3
rk1078 n643__chipdriverout n644__chipdriverout 226.6e-3
rk1079 n644__chipdriverout n645__chipdriverout 116.5e-3
rk1080 n645__chipdriverout n646__chipdriverout 365.7e-3
rk1081 n646__chipdriverout n647__chipdriverout 242.8e-3
rk1082 n647__chipdriverout n648__chipdriverout 119.7e-3
rk1084 n640__chipdriverout n641__chipdriverout 5.7692
rk1085 n640__chipdriverout n644__chipdriverout 3.75
rk1086 n640__chipdriverout n647__chipdriverout 3.75
rk1090 n6__x3 n3__x3 4.923e-3
rk1092 n6__y3 n3__y3 4.923e-3
rk1094 n368__vddio n383__vddio 30.13e-3
rk1095 n383__vddio n369__vddio 335.6e-3
rk1096 n369__vddio n372__vddio 343.1e-3
rk1097 n372__vddio n384__vddio 42.68e-3
rk1098 n384__vddio n373__vddio 321.2e-3
rk1099 n373__vddio n376__vddio 362.5e-3
rk1100 n376__vddio n385__vddio 40.17e-3
rk1101 n385__vddio n377__vddio 323.7e-3
rk1102 n377__vddio n380__vddio 343.1e-3
rk1103 n380__vddio n386__vddio 52.73e-3
rk1104 n386__vddio n387__vddio 394.2e-3
rk1105 n382__vddio n383__vddio 3.1
rk1106 n382__vddio n384__vddio 3.1
rk1107 n382__vddio n385__vddio 3.1
rk1108 n382__vddio n386__vddio 3.1
rk1109 n218__vss n215__vss 55.24e-3
rk1110 n215__vss n214__vss 365.7e-3
rk1111 n214__vss n219__vss 298.6e-3
rk1112 n219__vss n211__vss 42.68e-3
rk1113 n211__vss n210__vss 365.7e-3
rk1114 n210__vss n220__vss 187.7e-3
rk1115 n220__vss n221__vss 264.6e-3
rk1116 n217__vss n218__vss 3.75
rk1117 n217__vss n219__vss 3.75
rk1118 n217__vss n220__vss 5.7692
rk1119 n210__i1__i14__net1 n321__i1__i14__net1 125e-3
rk1120 n212__i1__i14__net1 n322__i1__i14__net1 125e-3
rk1122 n664__chipdriverout n666__chipdriverout 210.4e-3
rk1123 n666__chipdriverout n667__chipdriverout 155.3e-3
rk1124 n667__chipdriverout n668__chipdriverout 343.1e-3
rk1125 n668__chipdriverout n669__chipdriverout 226.6e-3
rk1126 n669__chipdriverout n670__chipdriverout 139.1e-3
rk1127 n670__chipdriverout n671__chipdriverout 362.5e-3
rk1128 n671__chipdriverout n672__chipdriverout 223.4e-3
rk1129 n672__chipdriverout n673__chipdriverout 142.4e-3
rk1130 n673__chipdriverout n674__chipdriverout 343.1e-3
rk1131 n674__chipdriverout n675__chipdriverout 239.6e-3
rk1132 n675__chipdriverout n676__chipdriverout 126.2e-3
rk1134 n665__chipdriverout n666__chipdriverout 3.1
rk1135 n665__chipdriverout n669__chipdriverout 3.1
rk1136 n665__chipdriverout n672__chipdriverout 3.1
rk1137 n665__chipdriverout n675__chipdriverout 3.1
rk1139 n680__chipdriverout n681__chipdriverout 12.55e-3
rk1140 n681__chipdriverout n682__chipdriverout 365.7e-3
rk1141 n682__chipdriverout n683__chipdriverout 226.6e-3
rk1142 n683__chipdriverout n684__chipdriverout 116.5e-3
rk1143 n684__chipdriverout n685__chipdriverout 365.7e-3
rk1144 n685__chipdriverout n686__chipdriverout 242.8e-3
rk1145 n686__chipdriverout n687__chipdriverout 119.7e-3
rk1147 n679__chipdriverout n680__chipdriverout 5.7692
rk1148 n679__chipdriverout n683__chipdriverout 3.75
rk1149 n679__chipdriverout n686__chipdriverout 3.75
rk1150 i5__i7__i0__i2__net21 n2__i5__i7__i0__i2__net21 62.1844
rk1151 i5__i7__i0__i2__net23 n2__i5__i7__i0__i2__net23 150.195
rk1152 i5__i7__i1__i2__net21 n2__i5__i7__i1__i2__net21 62.1844
rk1153 i5__i7__i1__i2__net23 n2__i5__i7__i1__i2__net23 150.195
rk1154 n218__i1__i14__net1 n329__i1__i14__net1 125e-3
rk1155 n220__i1__i14__net1 n330__i1__i14__net1 125e-3
rk1156 n64__i5__clk4 n47__i5__clk4 505.3e-3
rk1157 n30__i5__i7__i0__net1 n22__i5__i7__i0__net1 505.3e-3
rk1158 n68__i5__clk4 n49__i5__clk4 505.3e-3
rk1159 n30__i5__i7__i1__net1 n22__i5__i7__i1__net1 505.3e-3
rk1161 n388__vddio n404__vddio 30.13e-3
rk1162 n404__vddio n391__vddio 335.6e-3
rk1163 n391__vddio n392__vddio 343.1e-3
rk1164 n392__vddio n405__vddio 42.68e-3
rk1165 n405__vddio n395__vddio 321.2e-3
rk1166 n395__vddio n396__vddio 362.5e-3
rk1167 n396__vddio n406__vddio 40.17e-3
rk1168 n406__vddio n399__vddio 323.7e-3
rk1169 n399__vddio n400__vddio 343.1e-3
rk1170 n400__vddio n407__vddio 52.73e-3
rk1171 n407__vddio n408__vddio 394.2e-3
rk1172 n403__vddio n404__vddio 3.1
rk1173 n403__vddio n405__vddio 3.1
rk1174 n403__vddio n406__vddio 3.1
rk1175 n403__vddio n407__vddio 3.1
rk1176 n231__vss n229__vss 55.24e-3
rk1177 n229__vss n226__vss 365.7e-3
rk1178 n226__vss n232__vss 298.6e-3
rk1179 n232__vss n225__vss 42.68e-3
rk1180 n225__vss n222__vss 365.7e-3
rk1181 n222__vss n233__vss 187.7e-3
rk1182 n233__vss n234__vss 264.6e-3
rk1183 n230__vss n231__vss 3.75
rk1184 n230__vss n232__vss 3.75
rk1185 n230__vss n233__vss 5.7692
rk1186 n226__i1__i14__net1 n337__i1__i14__net1 125e-3
rk1187 n228__i1__i14__net1 n338__i1__i14__net1 125e-3
rk1189 n703__chipdriverout n705__chipdriverout 210.4e-3
rk1190 n705__chipdriverout n706__chipdriverout 155.3e-3
rk1191 n706__chipdriverout n707__chipdriverout 343.1e-3
rk1192 n707__chipdriverout n708__chipdriverout 226.6e-3
rk1193 n708__chipdriverout n709__chipdriverout 139.1e-3
rk1194 n709__chipdriverout n710__chipdriverout 362.5e-3
rk1195 n710__chipdriverout n711__chipdriverout 223.4e-3
rk1196 n711__chipdriverout n712__chipdriverout 142.4e-3
rk1197 n712__chipdriverout n713__chipdriverout 343.1e-3
rk1198 n713__chipdriverout n714__chipdriverout 239.6e-3
rk1199 n714__chipdriverout n715__chipdriverout 126.2e-3
rk1201 n704__chipdriverout n705__chipdriverout 3.1
rk1202 n704__chipdriverout n708__chipdriverout 3.1
rk1203 n704__chipdriverout n711__chipdriverout 3.1
rk1204 n704__chipdriverout n714__chipdriverout 3.1
rk1206 n719__chipdriverout n720__chipdriverout 12.55e-3
rk1207 n720__chipdriverout n721__chipdriverout 365.7e-3
rk1208 n721__chipdriverout n722__chipdriverout 226.6e-3
rk1209 n722__chipdriverout n723__chipdriverout 116.5e-3
rk1210 n723__chipdriverout n724__chipdriverout 365.7e-3
rk1211 n724__chipdriverout n725__chipdriverout 242.8e-3
rk1212 n725__chipdriverout n726__chipdriverout 119.7e-3
rk1214 n718__chipdriverout n719__chipdriverout 5.7692
rk1215 n718__chipdriverout n722__chipdriverout 3.75
rk1216 n718__chipdriverout n725__chipdriverout 3.75
rk1217 n5__i5__i7__i0__i2__net22 n6__i5__i7__i0__i2__net22 31.2679
rk1218 n6__i5__i7__i0__i2__net22 n7__i5__i7__i0__i2__net22 75.2632
rk1219 n6__i5__i7__i0__i2__net22 n3__i5__i7__i0__i2__net22 230.1e-3
rk1220 n5__i5__i7__i1__i2__net22 n6__i5__i7__i1__i2__net22 31.2679
rk1221 n6__i5__i7__i1__i2__net22 n7__i5__i7__i1__i2__net22 75.2632
rk1222 n6__i5__i7__i1__i2__net22 n3__i5__i7__i1__i2__net22 230.1e-3
rk1223 n238__i1__i14__net1 n349__i1__i14__net1 125e-3
rk1224 n240__i1__i14__net1 n350__i1__i14__net1 125e-3
rk1226 n409__vddio n429__vddio 30.13e-3
rk1227 n429__vddio n412__vddio 335.6e-3
rk1228 n412__vddio n413__vddio 343.1e-3
rk1229 n413__vddio n430__vddio 42.68e-3
rk1230 n430__vddio n416__vddio 321.2e-3
rk1231 n416__vddio n417__vddio 362.5e-3
rk1232 n417__vddio n431__vddio 40.17e-3
rk1233 n431__vddio n420__vddio 323.7e-3
rk1234 n420__vddio n421__vddio 343.1e-3
rk1235 n421__vddio n432__vddio 52.73e-3
rk1236 n432__vddio n433__vddio 394.2e-3
rk1237 n428__vddio n429__vddio 3.1
rk1238 n428__vddio n430__vddio 3.1
rk1239 n428__vddio n431__vddio 3.1
rk1240 n428__vddio n432__vddio 3.1
rk1241 n244__vss n242__vss 55.24e-3
rk1242 n242__vss n239__vss 365.7e-3
rk1243 n239__vss n245__vss 298.6e-3
rk1244 n245__vss n238__vss 42.68e-3
rk1245 n238__vss n235__vss 365.7e-3
rk1246 n235__vss n246__vss 187.7e-3
rk1247 n246__vss n247__vss 264.6e-3
rk1248 n243__vss n244__vss 3.75
rk1249 n243__vss n245__vss 3.75
rk1250 n243__vss n246__vss 5.7692
rk1251 n242__i1__i14__net1 n353__i1__i14__net1 125e-3
rk1252 n244__i1__i14__net1 n354__i1__i14__net1 125e-3
rk1253 i5__i7__i0__i2__net24 n2__i5__i7__i0__i2__net24 62.1844
rk1254 i5__i7__i0__i2__net25 n2__i5__i7__i0__i2__net25 150.195
rk1255 i5__i7__i1__i2__net24 n2__i5__i7__i1__i2__net24 62.1844
rk1256 i5__i7__i1__i2__net25 n2__i5__i7__i1__i2__net25 150.195
rk1257 n55__i5__clk4 n74__i5__clk4 4.923e-3
rk1258 n32__i5__i7__i0__net1 n26__i5__i7__i0__net1 507.7e-3
rk1259 n57__i5__clk4 n75__i5__clk4 4.923e-3
rk1260 n32__i5__i7__i1__net1 n26__i5__i7__i1__net1 507.7e-3
rk1262 n742__chipdriverout n744__chipdriverout 210.4e-3
rk1263 n744__chipdriverout n745__chipdriverout 155.3e-3
rk1264 n745__chipdriverout n746__chipdriverout 343.1e-3
rk1265 n746__chipdriverout n747__chipdriverout 226.6e-3
rk1266 n747__chipdriverout n748__chipdriverout 139.1e-3
rk1267 n748__chipdriverout n749__chipdriverout 362.5e-3
rk1268 n749__chipdriverout n750__chipdriverout 223.4e-3
rk1269 n750__chipdriverout n751__chipdriverout 142.4e-3
rk1270 n751__chipdriverout n752__chipdriverout 343.1e-3
rk1271 n752__chipdriverout n753__chipdriverout 239.6e-3
rk1272 n753__chipdriverout n754__chipdriverout 126.2e-3
rk1274 n743__chipdriverout n744__chipdriverout 3.1
rk1275 n743__chipdriverout n747__chipdriverout 3.1
rk1276 n743__chipdriverout n750__chipdriverout 3.1
rk1277 n743__chipdriverout n753__chipdriverout 3.1
rk1279 n758__chipdriverout n759__chipdriverout 12.55e-3
rk1280 n759__chipdriverout n760__chipdriverout 365.7e-3
rk1281 n760__chipdriverout n761__chipdriverout 226.6e-3
rk1282 n761__chipdriverout n762__chipdriverout 116.5e-3
rk1283 n762__chipdriverout n763__chipdriverout 365.7e-3
rk1284 n763__chipdriverout n764__chipdriverout 242.8e-3
rk1285 n764__chipdriverout n765__chipdriverout 119.7e-3
rk1287 n757__chipdriverout n758__chipdriverout 5.7692
rk1288 n757__chipdriverout n761__chipdriverout 3.75
rk1289 n757__chipdriverout n764__chipdriverout 3.75
rk1290 n254__i1__i14__net1 n365__i1__i14__net1 125e-3
rk1291 n256__i1__i14__net1 n366__i1__i14__net1 125e-3
rk1293 n435__vddio n450__vddio 30.13e-3
rk1294 n450__vddio n436__vddio 335.6e-3
rk1295 n436__vddio n439__vddio 343.1e-3
rk1296 n439__vddio n451__vddio 42.68e-3
rk1297 n451__vddio n440__vddio 321.2e-3
rk1298 n440__vddio n443__vddio 362.5e-3
rk1299 n443__vddio n452__vddio 40.17e-3
rk1300 n452__vddio n444__vddio 323.7e-3
rk1301 n444__vddio n447__vddio 343.1e-3
rk1302 n447__vddio n453__vddio 52.73e-3
rk1303 n453__vddio n454__vddio 394.2e-3
rk1304 n449__vddio n450__vddio 3.1
rk1305 n449__vddio n451__vddio 3.1
rk1306 n449__vddio n452__vddio 3.1
rk1307 n449__vddio n453__vddio 3.1
rk1308 n257__vss n254__vss 55.24e-3
rk1309 n254__vss n253__vss 365.7e-3
rk1310 n253__vss n258__vss 298.6e-3
rk1311 n258__vss n250__vss 42.68e-3
rk1312 n250__vss n249__vss 365.7e-3
rk1313 n249__vss n259__vss 187.7e-3
rk1314 n259__vss n260__vss 266.4e-3
rk1315 n256__vss n257__vss 3.75
rk1316 n256__vss n258__vss 3.75
rk1317 n256__vss n259__vss 5.7692
rk1318 n258__i1__i14__net1 n369__i1__i14__net1 125e-3
rk1319 n260__i1__i14__net1 n370__i1__i14__net1 125e-3
rk1320 n25__reset n32__reset 577.1e-3
rk1321 n27__reset n35__reset 77.13e-3
rk1323 n782__chipdriverout n783__chipdriverout 12.55e-3
rk1324 n783__chipdriverout n784__chipdriverout 365.7e-3
rk1325 n784__chipdriverout n785__chipdriverout 226.6e-3
rk1326 n785__chipdriverout n786__chipdriverout 116.5e-3
rk1327 n786__chipdriverout n787__chipdriverout 365.7e-3
rk1328 n787__chipdriverout n788__chipdriverout 242.8e-3
rk1329 n788__chipdriverout n789__chipdriverout 119.7e-3
rk1331 n781__chipdriverout n782__chipdriverout 5.7692
rk1332 n781__chipdriverout n785__chipdriverout 3.75
rk1333 n781__chipdriverout n788__chipdriverout 3.75
rk1335 n792__chipdriverout n794__chipdriverout 210.4e-3
rk1336 n794__chipdriverout n795__chipdriverout 155.3e-3
rk1337 n795__chipdriverout n796__chipdriverout 343.1e-3
rk1338 n796__chipdriverout n797__chipdriverout 226.6e-3
rk1339 n797__chipdriverout n798__chipdriverout 139.1e-3
rk1340 n798__chipdriverout n799__chipdriverout 362.5e-3
rk1341 n799__chipdriverout n800__chipdriverout 223.4e-3
rk1342 n800__chipdriverout n801__chipdriverout 142.4e-3
rk1343 n801__chipdriverout n802__chipdriverout 343.1e-3
rk1344 n802__chipdriverout n803__chipdriverout 239.6e-3
rk1345 n803__chipdriverout n804__chipdriverout 126.2e-3
rk1347 n793__chipdriverout n794__chipdriverout 3.1
rk1348 n793__chipdriverout n797__chipdriverout 3.1
rk1349 n793__chipdriverout n800__chipdriverout 3.1
rk1350 n793__chipdriverout n803__chipdriverout 3.1
rk1351 n4__i5__i7__x3out n5__i5__i7__x3out 19.2986
rk1352 n5__i5__i7__x3out n7__i5__i7__x3out 528.7e-3
rk1353 n7__i5__i7__x3out n8__i5__i7__x3out 75.4978
rk1354 n6__i5__i7__x3out n7__i5__i7__x3out 31
rk1355 n6__i5__i7__y3out n7__i5__i7__y3out 19.2986
rk1356 n7__i5__i7__y3out n9__i5__i7__y3out 528.7e-3
rk1357 n9__i5__i7__y3out n10__i5__i7__y3out 75.4978
rk1358 n8__i5__i7__y3out n9__i5__i7__y3out 31
rk1359 n270__i1__i14__net1 n377__i1__i14__net1 125e-3
rk1360 n272__i1__i14__net1 n378__i1__i14__net1 125e-3
rk1362 n462__vddio n464__vddio 30.13e-3
rk1363 n464__vddio n465__vddio 335.6e-3
rk1364 n465__vddio n466__vddio 343.1e-3
rk1365 n466__vddio n467__vddio 42.68e-3
rk1366 n467__vddio n468__vddio 321.2e-3
rk1367 n468__vddio n469__vddio 362.5e-3
rk1368 n469__vddio n470__vddio 40.17e-3
rk1369 n470__vddio n471__vddio 323.7e-3
rk1370 n471__vddio n472__vddio 343.1e-3
rk1371 n472__vddio n473__vddio 52.73e-3
rk1372 n473__vddio n474__vddio 394.2e-3
rk1373 n463__vddio n464__vddio 3.1
rk1374 n463__vddio n467__vddio 3.1
rk1375 n463__vddio n470__vddio 3.1
rk1376 n463__vddio n473__vddio 3.1
rk1377 n262__vss n263__vss 55.24e-3
rk1378 n263__vss n264__vss 365.7e-3
rk1379 n264__vss n265__vss 298.6e-3
rk1380 n265__vss n266__vss 42.68e-3
rk1381 n266__vss n267__vss 365.7e-3
rk1382 n267__vss n268__vss 187.7e-3
rk1383 n268__vss n269__vss 264.6e-3
rk1384 n261__vss n262__vss 3.75
rk1385 n261__vss n265__vss 3.75
rk1386 n261__vss n268__vss 5.7692
rk1387 n274__i1__i14__net1 n385__i1__i14__net1 125e-3
rk1388 n276__i1__i14__net1 n386__i1__i14__net1 125e-3
rk1389 n2__i5__i7__y2out n14__i5__i7__y2out 45.2869
rk1390 n9__i5__i7__y1out n13__i5__i7__y1out 45.2869
rk1392 n821__chipdriverout n822__chipdriverout 12.55e-3
rk1393 n822__chipdriverout n823__chipdriverout 365.7e-3
rk1394 n823__chipdriverout n824__chipdriverout 226.6e-3
rk1395 n824__chipdriverout n825__chipdriverout 116.5e-3
rk1396 n825__chipdriverout n826__chipdriverout 365.7e-3
rk1397 n826__chipdriverout n827__chipdriverout 242.8e-3
rk1398 n827__chipdriverout n828__chipdriverout 119.7e-3
rk1400 n820__chipdriverout n821__chipdriverout 5.7692
rk1401 n820__chipdriverout n824__chipdriverout 3.75
rk1402 n820__chipdriverout n827__chipdriverout 3.75
rk1404 n831__chipdriverout n833__chipdriverout 210.4e-3
rk1405 n833__chipdriverout n834__chipdriverout 155.3e-3
rk1406 n834__chipdriverout n835__chipdriverout 343.1e-3
rk1407 n835__chipdriverout n836__chipdriverout 226.6e-3
rk1408 n836__chipdriverout n837__chipdriverout 139.1e-3
rk1409 n837__chipdriverout n838__chipdriverout 362.5e-3
rk1410 n838__chipdriverout n839__chipdriverout 223.4e-3
rk1411 n839__chipdriverout n840__chipdriverout 142.4e-3
rk1412 n840__chipdriverout n841__chipdriverout 343.1e-3
rk1413 n841__chipdriverout n842__chipdriverout 239.6e-3
rk1414 n842__chipdriverout n843__chipdriverout 126.2e-3
rk1416 n832__chipdriverout n833__chipdriverout 3.1
rk1417 n832__chipdriverout n836__chipdriverout 3.1
rk1418 n832__chipdriverout n839__chipdriverout 3.1
rk1419 n832__chipdriverout n842__chipdriverout 3.1
rk1423 n483__vddio n485__vddio 30.13e-3
rk1424 n485__vddio n486__vddio 335.6e-3
rk1425 n486__vddio n487__vddio 343.1e-3
rk1426 n487__vddio n488__vddio 42.68e-3
rk1427 n488__vddio n489__vddio 321.2e-3
rk1428 n489__vddio n490__vddio 362.5e-3
rk1429 n490__vddio n491__vddio 40.17e-3
rk1430 n491__vddio n492__vddio 323.7e-3
rk1431 n492__vddio n493__vddio 343.1e-3
rk1432 n493__vddio n494__vddio 52.73e-3
rk1433 n494__vddio n495__vddio 394.2e-3
rk1434 n484__vddio n485__vddio 3.1
rk1435 n484__vddio n488__vddio 3.1
rk1436 n484__vddio n491__vddio 3.1
rk1437 n484__vddio n494__vddio 3.1
rk1438 n275__vss n276__vss 55.24e-3
rk1439 n276__vss n277__vss 365.7e-3
rk1440 n277__vss n278__vss 298.6e-3
rk1441 n278__vss n279__vss 42.68e-3
rk1442 n279__vss n280__vss 365.7e-3
rk1443 n280__vss n281__vss 187.7e-3
rk1444 n281__vss n282__vss 264.6e-3
rk1445 n274__vss n275__vss 3.75
rk1446 n274__vss n278__vss 3.75
rk1447 n274__vss n281__vss 5.7692
rk1448 n294__i1__i14__net1 n401__i1__i14__net1 125e-3
rk1449 n296__i1__i14__net1 n402__i1__i14__net1 125e-3
rk1451 n859__chipdriverout n861__chipdriverout 210.4e-3
rk1452 n861__chipdriverout n862__chipdriverout 155.3e-3
rk1453 n862__chipdriverout n863__chipdriverout 343.1e-3
rk1454 n863__chipdriverout n864__chipdriverout 226.6e-3
rk1455 n864__chipdriverout n865__chipdriverout 139.1e-3
rk1456 n865__chipdriverout n866__chipdriverout 362.5e-3
rk1457 n866__chipdriverout n867__chipdriverout 223.4e-3
rk1458 n867__chipdriverout n868__chipdriverout 142.4e-3
rk1459 n868__chipdriverout n869__chipdriverout 343.1e-3
rk1460 n869__chipdriverout n870__chipdriverout 239.6e-3
rk1461 n870__chipdriverout n871__chipdriverout 126.2e-3
rk1463 n860__chipdriverout n861__chipdriverout 3.1
rk1464 n860__chipdriverout n864__chipdriverout 3.1
rk1465 n860__chipdriverout n867__chipdriverout 3.1
rk1466 n860__chipdriverout n870__chipdriverout 3.1
rk1468 n883__chipdriverout n884__chipdriverout 12.55e-3
rk1469 n884__chipdriverout n885__chipdriverout 365.7e-3
rk1470 n885__chipdriverout n886__chipdriverout 226.6e-3
rk1471 n886__chipdriverout n887__chipdriverout 116.5e-3
rk1472 n887__chipdriverout n888__chipdriverout 365.7e-3
rk1473 n888__chipdriverout n889__chipdriverout 242.8e-3
rk1474 n889__chipdriverout n890__chipdriverout 119.7e-3
rk1476 n882__chipdriverout n883__chipdriverout 5.7692
rk1477 n882__chipdriverout n886__chipdriverout 3.75
rk1478 n882__chipdriverout n889__chipdriverout 3.75
rk1479 n302__i1__i14__net1 n409__i1__i14__net1 125e-3
rk1480 n304__i1__i14__net1 n410__i1__i14__net1 125e-3
rk1482 n504__vddio n506__vddio 30.13e-3
rk1483 n506__vddio n507__vddio 335.6e-3
rk1484 n507__vddio n508__vddio 343.1e-3
rk1485 n508__vddio n509__vddio 42.68e-3
rk1486 n509__vddio n510__vddio 321.2e-3
rk1487 n510__vddio n511__vddio 362.5e-3
rk1488 n511__vddio n512__vddio 40.17e-3
rk1489 n512__vddio n513__vddio 323.7e-3
rk1490 n513__vddio n514__vddio 343.1e-3
rk1491 n514__vddio n515__vddio 52.73e-3
rk1492 n515__vddio n516__vddio 394.2e-3
rk1493 n505__vddio n506__vddio 3.1
rk1494 n505__vddio n509__vddio 3.1
rk1495 n505__vddio n512__vddio 3.1
rk1496 n505__vddio n515__vddio 3.1
rk1497 n292__vss n289__vss 55.24e-3
rk1498 n289__vss n288__vss 365.7e-3
rk1499 n288__vss n293__vss 298.6e-3
rk1500 n293__vss n294__vss 42.68e-3
rk1501 n294__vss n295__vss 365.7e-3
rk1502 n295__vss n296__vss 187.7e-3
rk1503 n296__vss n297__vss 264.6e-3
rk1504 n291__vss n292__vss 3.75
rk1505 n291__vss n293__vss 3.75
rk1506 n291__vss n296__vss 5.7692
rk1507 n5__i5__i7__xor2 n6__i5__i7__xor2 33.29e-3
rk1508 n6__i5__i7__xor2 n4__i5__i7__xor2 31.0291
rk1509 n4__i5__i7__xor2 n5__i5__i7__xor2 31
rk1510 n7__i5__i7__xor2 n8__i5__i7__xor2 75.0296
rk1511 n8__i5__i7__xor2 n7__i5__i7__xor2 75.0338
rk1512 n5__i5__i7__xor1 n6__i5__i7__xor1 33.29e-3
rk1513 n6__i5__i7__xor1 n4__i5__i7__xor1 31.0291
rk1514 n4__i5__i7__xor1 n5__i5__i7__xor1 31
rk1515 n7__i5__i7__xor1 n8__i5__i7__xor1 75.0296
rk1516 n8__i5__i7__xor1 n7__i5__i7__xor1 75.0338
rk1517 n305__i1__i14__net1 n417__i1__i14__net1 125e-3
rk1518 n307__i1__i14__net1 n418__i1__i14__net1 125e-3
rk1519 n3__i5__i7__i8__net1 n5__i5__i7__i8__net1 31.3722
rk1520 n5__i5__i7__i8__net1 n7__i5__i7__i8__net1 204.7e-3
rk1521 n7__i5__i7__i8__net1 n2__i5__i7__i8__net1 399.2e-3
rk1522 n4__i5__i7__i8__net1 n5__i5__i7__i8__net1 75
rk1523 n6__i5__i7__i8__net1 n7__i5__i7__i8__net1 75
rk1524 n3__i5__i7__i3__net1 n5__i5__i7__i3__net1 31.3722
rk1525 n5__i5__i7__i3__net1 n7__i5__i7__i3__net1 204.7e-3
rk1526 n7__i5__i7__i3__net1 n2__i5__i7__i3__net1 399.2e-3
rk1527 n4__i5__i7__i3__net1 n5__i5__i7__i3__net1 75
rk1528 n6__i5__i7__i3__net1 n7__i5__i7__i3__net1 75
rk1529 n12__i5__i7__y2out n16__i5__i7__y2out 292e-3
rk1530 n16__i5__i7__y2out n17__i5__i7__y2out 31.1232
rk1531 n12__i5__i7__y1out n16__i5__i7__y1out 292e-3
rk1532 n16__i5__i7__y1out n17__i5__i7__y1out 31.1232
rk1534 n899__chipdriverout n900__chipdriverout 12.55e-3
rk1535 n900__chipdriverout n901__chipdriverout 365.7e-3
rk1536 n901__chipdriverout n902__chipdriverout 226.6e-3
rk1537 n902__chipdriverout n903__chipdriverout 116.5e-3
rk1538 n903__chipdriverout n904__chipdriverout 365.7e-3
rk1539 n904__chipdriverout n905__chipdriverout 242.8e-3
rk1540 n905__chipdriverout n906__chipdriverout 119.7e-3
rk1542 n898__chipdriverout n899__chipdriverout 5.7692
rk1543 n898__chipdriverout n902__chipdriverout 3.75
rk1544 n898__chipdriverout n905__chipdriverout 3.75
rk1546 n909__chipdriverout n911__chipdriverout 210.4e-3
rk1547 n911__chipdriverout n912__chipdriverout 155.3e-3
rk1548 n912__chipdriverout n913__chipdriverout 343.1e-3
rk1549 n913__chipdriverout n914__chipdriverout 226.6e-3
rk1550 n914__chipdriverout n915__chipdriverout 139.1e-3
rk1551 n915__chipdriverout n916__chipdriverout 362.5e-3
rk1552 n916__chipdriverout n917__chipdriverout 223.4e-3
rk1553 n917__chipdriverout n918__chipdriverout 142.4e-3
rk1554 n918__chipdriverout n919__chipdriverout 343.1e-3
rk1555 n919__chipdriverout n920__chipdriverout 239.6e-3
rk1556 n920__chipdriverout n921__chipdriverout 126.2e-3
rk1558 n910__chipdriverout n911__chipdriverout 3.1
rk1559 n910__chipdriverout n914__chipdriverout 3.1
rk1560 n910__chipdriverout n917__chipdriverout 3.1
rk1561 n910__chipdriverout n920__chipdriverout 3.1
rk1562 n14__i5__i7__x2out n15__i5__i7__x2out 31.115
rk1563 n15__i5__i7__x2out n16__i5__i7__x2out 328.8e-3
rk1564 n16__i5__i7__x2out n13__i5__i7__x2out 11.8e-3
rk1565 n15__i5__i7__x2out n17__i5__i7__x2out 75.115
rk1566 n2__i5__i7__x2out n16__i5__i7__x2out 15
rk1567 n14__i5__i7__x1out n15__i5__i7__x1out 31.115
rk1568 n15__i5__i7__x1out n16__i5__i7__x1out 328.8e-3
rk1569 n16__i5__i7__x1out n13__i5__i7__x1out 11.8e-3
rk1570 n15__i5__i7__x1out n17__i5__i7__x1out 75.115
rk1571 n9__i5__i7__x1out n16__i5__i7__x1out 15
rk1575 n525__vddio n527__vddio 30.13e-3
rk1576 n527__vddio n528__vddio 335.6e-3
rk1577 n528__vddio n529__vddio 343.1e-3
rk1578 n529__vddio n530__vddio 42.68e-3
rk1579 n530__vddio n531__vddio 321.2e-3
rk1580 n531__vddio n532__vddio 362.5e-3
rk1581 n532__vddio n533__vddio 40.17e-3
rk1582 n533__vddio n534__vddio 323.7e-3
rk1583 n534__vddio n535__vddio 343.1e-3
rk1584 n535__vddio n536__vddio 52.73e-3
rk1585 n536__vddio n537__vddio 394.2e-3
rk1586 n526__vddio n527__vddio 3.1
rk1587 n526__vddio n530__vddio 3.1
rk1588 n526__vddio n533__vddio 3.1
rk1589 n526__vddio n536__vddio 3.1
rk1590 n309__vss n306__vss 55.24e-3
rk1591 n306__vss n305__vss 369.4e-3
rk1592 n305__vss n310__vss 304e-3
rk1593 n310__vss n302__vss 42.68e-3
rk1594 n302__vss n301__vss 369.4e-3
rk1595 n301__vss n311__vss 189.5e-3
rk1596 n311__vss n312__vss 264.6e-3
rk1597 n308__vss n309__vss 3.75
rk1598 n308__vss n310__vss 3.75
rk1599 n308__vss n311__vss 5.7692
rk1600 n325__i1__i14__net1 n437__i1__i14__net1 125e-3
rk1601 n327__i1__i14__net1 n438__i1__i14__net1 125e-3
rk1603 n938__chipdriverout n939__chipdriverout 12.55e-3
rk1604 n939__chipdriverout n940__chipdriverout 365.7e-3
rk1605 n940__chipdriverout n941__chipdriverout 226.6e-3
rk1606 n941__chipdriverout n942__chipdriverout 116.5e-3
rk1607 n942__chipdriverout n943__chipdriverout 365.7e-3
rk1608 n943__chipdriverout n944__chipdriverout 242.8e-3
rk1609 n944__chipdriverout n945__chipdriverout 119.7e-3
rk1611 n937__chipdriverout n938__chipdriverout 5.7692
rk1612 n937__chipdriverout n941__chipdriverout 3.75
rk1613 n937__chipdriverout n944__chipdriverout 3.75
rk1615 n948__chipdriverout n950__chipdriverout 210.4e-3
rk1616 n950__chipdriverout n951__chipdriverout 155.3e-3
rk1617 n951__chipdriverout n952__chipdriverout 343.1e-3
rk1618 n952__chipdriverout n953__chipdriverout 226.6e-3
rk1619 n953__chipdriverout n954__chipdriverout 139.1e-3
rk1620 n954__chipdriverout n955__chipdriverout 362.5e-3
rk1621 n955__chipdriverout n956__chipdriverout 223.4e-3
rk1622 n956__chipdriverout n957__chipdriverout 142.4e-3
rk1623 n957__chipdriverout n958__chipdriverout 343.1e-3
rk1624 n958__chipdriverout n959__chipdriverout 239.6e-3
rk1625 n959__chipdriverout n960__chipdriverout 126.2e-3
rk1627 n949__chipdriverout n950__chipdriverout 3.1
rk1628 n949__chipdriverout n953__chipdriverout 3.1
rk1629 n949__chipdriverout n956__chipdriverout 3.1
rk1630 n949__chipdriverout n959__chipdriverout 3.1
rk1634 n546__vddio n561__vddio 30.13e-3
rk1635 n561__vddio n547__vddio 335.6e-3
rk1636 n547__vddio n550__vddio 343.1e-3
rk1637 n550__vddio n562__vddio 42.68e-3
rk1638 n562__vddio n551__vddio 321.2e-3
rk1639 n551__vddio n554__vddio 362.5e-3
rk1640 n554__vddio n563__vddio 40.17e-3
rk1641 n563__vddio n555__vddio 323.7e-3
rk1642 n555__vddio n558__vddio 343.1e-3
rk1643 n558__vddio n564__vddio 52.73e-3
rk1644 n564__vddio n565__vddio 394.2e-3
rk1645 n560__vddio n561__vddio 3.1
rk1646 n560__vddio n562__vddio 3.1
rk1647 n560__vddio n563__vddio 3.1
rk1648 n560__vddio n564__vddio 3.1
rk1649 n322__vss n319__vss 55.24e-3
rk1650 n319__vss n318__vss 365.7e-3
rk1651 n318__vss n323__vss 298.6e-3
rk1652 n323__vss n315__vss 42.68e-3
rk1653 n315__vss n314__vss 365.7e-3
rk1654 n314__vss n324__vss 187.7e-3
rk1655 n324__vss n325__vss 264.6e-3
rk1656 n321__vss n322__vss 3.75
rk1657 n321__vss n323__vss 3.75
rk1658 n321__vss n324__vss 5.7692
rk1659 n2__i5__i7__y3out n12__i5__i7__y3out 45.2869
rk1660 n9__i5__i7__y0out n13__i5__i7__y0out 45.2869
rk1661 n341__i1__i14__net1 n453__i1__i14__net1 125e-3
rk1662 n343__i1__i14__net1 n454__i1__i14__net1 125e-3
rk1664 n1003__chipdriverout n976__chipdriverout 12.55e-3
rk1665 n976__chipdriverout n977__chipdriverout 365.7e-3
rk1666 n977__chipdriverout n1004__chipdriverout 226.6e-3
rk1667 n1004__chipdriverout n980__chipdriverout 116.5e-3
rk1668 n980__chipdriverout n981__chipdriverout 365.7e-3
rk1669 n981__chipdriverout n1005__chipdriverout 242.8e-3
rk1670 n1005__chipdriverout n984__chipdriverout 119.7e-3
rk1672 n1002__chipdriverout n1003__chipdriverout 5.7692
rk1673 n1002__chipdriverout n1004__chipdriverout 3.75
rk1674 n1002__chipdriverout n1005__chipdriverout 3.75
rk1676 n985__chipdriverout n1009__chipdriverout 210.4e-3
rk1677 n1009__chipdriverout n988__chipdriverout 155.3e-3
rk1678 n988__chipdriverout n989__chipdriverout 343.1e-3
rk1679 n989__chipdriverout n1010__chipdriverout 226.6e-3
rk1680 n1010__chipdriverout n992__chipdriverout 139.1e-3
rk1681 n992__chipdriverout n993__chipdriverout 362.5e-3
rk1682 n993__chipdriverout n1011__chipdriverout 223.4e-3
rk1683 n1011__chipdriverout n996__chipdriverout 142.4e-3
rk1684 n996__chipdriverout n997__chipdriverout 343.1e-3
rk1685 n997__chipdriverout n1012__chipdriverout 239.6e-3
rk1686 n1012__chipdriverout n1000__chipdriverout 126.2e-3
rk1688 n1008__chipdriverout n1009__chipdriverout 3.1
rk1689 n1008__chipdriverout n1010__chipdriverout 3.1
rk1690 n1008__chipdriverout n1011__chipdriverout 3.1
rk1691 n1008__chipdriverout n1012__chipdriverout 3.1
rk1692 n346__i1__i14__net1 n461__i1__i14__net1 125e-3
rk1693 n348__i1__i14__net1 n462__i1__i14__net1 125e-3
rk1695 n577__vddio n579__vddio 30.13e-3
rk1696 n579__vddio n580__vddio 335.6e-3
rk1697 n580__vddio n581__vddio 343.1e-3
rk1698 n581__vddio n582__vddio 42.68e-3
rk1699 n582__vddio n583__vddio 321.2e-3
rk1700 n583__vddio n584__vddio 362.5e-3
rk1701 n584__vddio n585__vddio 40.17e-3
rk1702 n585__vddio n586__vddio 323.7e-3
rk1703 n586__vddio n587__vddio 343.1e-3
rk1704 n587__vddio n588__vddio 52.73e-3
rk1705 n588__vddio n589__vddio 394.2e-3
rk1706 n578__vddio n579__vddio 3.1
rk1707 n578__vddio n582__vddio 3.1
rk1708 n578__vddio n585__vddio 3.1
rk1709 n578__vddio n588__vddio 3.1
rk1710 n335__vss n332__vss 55.24e-3
rk1711 n332__vss n331__vss 369.4e-3
rk1712 n331__vss n336__vss 304e-3
rk1713 n336__vss n328__vss 42.68e-3
rk1714 n328__vss n327__vss 369.4e-3
rk1715 n327__vss n337__vss 189.5e-3
rk1716 n337__vss n338__vss 264.6e-3
rk1717 n334__vss n335__vss 3.75
rk1718 n334__vss n336__vss 3.75
rk1719 n334__vss n337__vss 5.7692
rk1723 n1016__chipdriverout n1017__chipdriverout 12.55e-3
rk1724 n1017__chipdriverout n1018__chipdriverout 365.7e-3
rk1725 n1018__chipdriverout n1019__chipdriverout 226.6e-3
rk1726 n1019__chipdriverout n1020__chipdriverout 116.5e-3
rk1727 n1020__chipdriverout n1021__chipdriverout 365.7e-3
rk1728 n1021__chipdriverout n1022__chipdriverout 242.8e-3
rk1729 n1022__chipdriverout n1023__chipdriverout 119.7e-3
rk1731 n1015__chipdriverout n1016__chipdriverout 5.7692
rk1732 n1015__chipdriverout n1019__chipdriverout 3.75
rk1733 n1015__chipdriverout n1022__chipdriverout 3.75
rk1735 n1026__chipdriverout n1028__chipdriverout 212.2e-3
rk1736 n1028__chipdriverout n1029__chipdriverout 157.2e-3
rk1737 n1029__chipdriverout n1030__chipdriverout 346.7e-3
rk1738 n1030__chipdriverout n1031__chipdriverout 228.4e-3
rk1739 n1031__chipdriverout n1032__chipdriverout 141e-3
rk1740 n1032__chipdriverout n1033__chipdriverout 366.1e-3
rk1741 n1033__chipdriverout n1034__chipdriverout 225.2e-3
rk1742 n1034__chipdriverout n1035__chipdriverout 144.2e-3
rk1743 n1035__chipdriverout n1036__chipdriverout 346.7e-3
rk1744 n1036__chipdriverout n1037__chipdriverout 241.4e-3
rk1745 n1037__chipdriverout n1038__chipdriverout 128e-3
rk1747 n1027__chipdriverout n1028__chipdriverout 3.1
rk1748 n1027__chipdriverout n1031__chipdriverout 3.1
rk1749 n1027__chipdriverout n1034__chipdriverout 3.1
rk1750 n1027__chipdriverout n1037__chipdriverout 3.1
rk1751 n362__i1__i14__net1 n473__i1__i14__net1 125e-3
rk1752 n364__i1__i14__net1 n474__i1__i14__net1 125e-3
rk1753 n5__i5__i7__xor3 n6__i5__i7__xor3 33.29e-3
rk1754 n6__i5__i7__xor3 n4__i5__i7__xor3 31.0291
rk1755 n4__i5__i7__xor3 n5__i5__i7__xor3 31
rk1756 n7__i5__i7__xor3 n8__i5__i7__xor3 75.0296
rk1757 n8__i5__i7__xor3 n7__i5__i7__xor3 75.0338
rk1758 n5__i5__i7__xor0 n6__i5__i7__xor0 33.29e-3
rk1759 n6__i5__i7__xor0 n4__i5__i7__xor0 31.0291
rk1760 n4__i5__i7__xor0 n5__i5__i7__xor0 31
rk1761 n7__i5__i7__xor0 n8__i5__i7__xor0 75.0296
rk1762 n8__i5__i7__xor0 n7__i5__i7__xor0 75.0338
rk1763 n348__vss n345__vss 55.24e-3
rk1764 n345__vss n344__vss 365.7e-3
rk1765 n344__vss n349__vss 298.6e-3
rk1766 n349__vss n341__vss 42.68e-3
rk1767 n341__vss n340__vss 365.7e-3
rk1768 n340__vss n350__vss 187.7e-3
rk1769 n350__vss n351__vss 264.6e-3
rk1770 n347__vss n348__vss 3.75
rk1771 n347__vss n349__vss 3.75
rk1772 n347__vss n350__vss 5.7692
rk1774 n598__vddio n613__vddio 30.13e-3
rk1775 n613__vddio n599__vddio 335.6e-3
rk1776 n599__vddio n602__vddio 343.1e-3
rk1777 n602__vddio n614__vddio 42.68e-3
rk1778 n614__vddio n603__vddio 321.2e-3
rk1779 n603__vddio n606__vddio 362.5e-3
rk1780 n606__vddio n615__vddio 40.17e-3
rk1781 n615__vddio n607__vddio 323.7e-3
rk1782 n607__vddio n610__vddio 343.1e-3
rk1783 n610__vddio n616__vddio 52.73e-3
rk1784 n616__vddio n617__vddio 394.2e-3
rk1785 n612__vddio n613__vddio 3.1
rk1786 n612__vddio n614__vddio 3.1
rk1787 n612__vddio n615__vddio 3.1
rk1788 n612__vddio n616__vddio 3.1
rk1789 n3__i5__i7__i9__net1 n5__i5__i7__i9__net1 31.3722
rk1790 n5__i5__i7__i9__net1 n7__i5__i7__i9__net1 204.7e-3
rk1791 n7__i5__i7__i9__net1 n2__i5__i7__i9__net1 399.2e-3
rk1792 n4__i5__i7__i9__net1 n5__i5__i7__i9__net1 75
rk1793 n6__i5__i7__i9__net1 n7__i5__i7__i9__net1 75
rk1794 n3__i5__i7__i2__net1 n5__i5__i7__i2__net1 31.3722
rk1795 n5__i5__i7__i2__net1 n7__i5__i7__i2__net1 204.7e-3
rk1796 n7__i5__i7__i2__net1 n2__i5__i7__i2__net1 399.2e-3
rk1797 n4__i5__i7__i2__net1 n5__i5__i7__i2__net1 75
rk1798 n6__i5__i7__i2__net1 n7__i5__i7__i2__net1 75
rk1799 n5__i5__i7__y3out n14__i5__i7__y3out 292e-3
rk1800 n14__i5__i7__y3out n15__i5__i7__y3out 31.1232
rk1801 n12__i5__i7__y0out n16__i5__i7__y0out 292e-3
rk1802 n16__i5__i7__y0out n17__i5__i7__y0out 31.1232
rk1803 n373__i1__i14__net1 n485__i1__i14__net1 125e-3
rk1804 n375__i1__i14__net1 n486__i1__i14__net1 125e-3
rk1805 n14__i5__i7__x3out n15__i5__i7__x3out 31.115
rk1806 n15__i5__i7__x3out n16__i5__i7__x3out 328.8e-3
rk1807 n16__i5__i7__x3out n13__i5__i7__x3out 11.8e-3
rk1808 n15__i5__i7__x3out n17__i5__i7__x3out 75.115
rk1809 n2__i5__i7__x3out n16__i5__i7__x3out 15
rk1810 n14__i5__i7__x0out n15__i5__i7__x0out 31.115
rk1811 n15__i5__i7__x0out n16__i5__i7__x0out 328.8e-3
rk1812 n16__i5__i7__x0out n13__i5__i7__x0out 11.8e-3
rk1813 n15__i5__i7__x0out n17__i5__i7__x0out 75.115
rk1814 n9__i5__i7__x0out n16__i5__i7__x0out 15
rk1816 n1055__chipdriverout n1056__chipdriverout 12.55e-3
rk1817 n1056__chipdriverout n1057__chipdriverout 365.7e-3
rk1818 n1057__chipdriverout n1058__chipdriverout 226.6e-3
rk1819 n1058__chipdriverout n1059__chipdriverout 116.5e-3
rk1820 n1059__chipdriverout n1060__chipdriverout 365.7e-3
rk1821 n1060__chipdriverout n1061__chipdriverout 242.8e-3
rk1822 n1061__chipdriverout n1062__chipdriverout 119.7e-3
rk1824 n1054__chipdriverout n1055__chipdriverout 5.7692
rk1825 n1054__chipdriverout n1058__chipdriverout 3.75
rk1826 n1054__chipdriverout n1061__chipdriverout 3.75
rk1828 n1065__chipdriverout n1067__chipdriverout 212.2e-3
rk1829 n1067__chipdriverout n1068__chipdriverout 157.2e-3
rk1830 n1068__chipdriverout n1069__chipdriverout 346.7e-3
rk1831 n1069__chipdriverout n1070__chipdriverout 228.4e-3
rk1832 n1070__chipdriverout n1071__chipdriverout 141e-3
rk1833 n1071__chipdriverout n1072__chipdriverout 366.1e-3
rk1834 n1072__chipdriverout n1073__chipdriverout 225.2e-3
rk1835 n1073__chipdriverout n1074__chipdriverout 144.2e-3
rk1836 n1074__chipdriverout n1075__chipdriverout 346.7e-3
rk1837 n1075__chipdriverout n1076__chipdriverout 241.4e-3
rk1838 n1076__chipdriverout n1077__chipdriverout 128e-3
rk1840 n1066__chipdriverout n1067__chipdriverout 3.1
rk1841 n1066__chipdriverout n1070__chipdriverout 3.1
rk1842 n1066__chipdriverout n1073__chipdriverout 3.1
rk1843 n1066__chipdriverout n1076__chipdriverout 3.1
rk1844 n380__i1__i14__net1 n489__i1__i14__net1 125e-3
rk1845 n382__i1__i14__net1 n490__i1__i14__net1 125e-3
rk1846 n353__vss n354__vss 55.24e-3
rk1847 n354__vss n355__vss 365.7e-3
rk1848 n355__vss n356__vss 298.6e-3
rk1849 n356__vss n357__vss 42.68e-3
rk1850 n357__vss n358__vss 365.7e-3
rk1851 n358__vss n359__vss 187.7e-3
rk1852 n359__vss n360__vss 264.6e-3
rk1853 n352__vss n353__vss 3.75
rk1854 n352__vss n356__vss 3.75
rk1855 n352__vss n359__vss 5.7692
rk1857 n619__vddio n621__vddio 30.13e-3
rk1858 n621__vddio n622__vddio 335.6e-3
rk1859 n622__vddio n623__vddio 343.1e-3
rk1860 n623__vddio n624__vddio 42.68e-3
rk1861 n624__vddio n625__vddio 321.2e-3
rk1862 n625__vddio n626__vddio 362.5e-3
rk1863 n626__vddio n627__vddio 40.17e-3
rk1864 n627__vddio n628__vddio 323.7e-3
rk1865 n628__vddio n629__vddio 343.1e-3
rk1866 n629__vddio n630__vddio 52.73e-3
rk1867 n630__vddio n631__vddio 394.2e-3
rk1868 n620__vddio n621__vddio 3.1
rk1869 n620__vddio n624__vddio 3.1
rk1870 n620__vddio n627__vddio 3.1
rk1871 n620__vddio n630__vddio 3.1
rk1872 n389__i1__i14__net1 n501__i1__i14__net1 125e-3
rk1873 n391__i1__i14__net1 n502__i1__i14__net1 125e-3
rk1875 n1120__chipdriverout n1093__chipdriverout 12.55e-3
rk1876 n1093__chipdriverout n1094__chipdriverout 365.7e-3
rk1877 n1094__chipdriverout n1121__chipdriverout 226.6e-3
rk1878 n1121__chipdriverout n1097__chipdriverout 116.5e-3
rk1879 n1097__chipdriverout n1098__chipdriverout 365.7e-3
rk1880 n1098__chipdriverout n1122__chipdriverout 242.8e-3
rk1881 n1122__chipdriverout n1101__chipdriverout 119.7e-3
rk1883 n1119__chipdriverout n1120__chipdriverout 5.7692
rk1884 n1119__chipdriverout n1121__chipdriverout 3.75
rk1885 n1119__chipdriverout n1122__chipdriverout 3.75
rk1887 n1102__chipdriverout n1126__chipdriverout 210.4e-3
rk1888 n1126__chipdriverout n1105__chipdriverout 155.3e-3
rk1889 n1105__chipdriverout n1106__chipdriverout 343.1e-3
rk1890 n1106__chipdriverout n1127__chipdriverout 226.6e-3
rk1891 n1127__chipdriverout n1109__chipdriverout 139.1e-3
rk1892 n1109__chipdriverout n1110__chipdriverout 362.5e-3
rk1893 n1110__chipdriverout n1128__chipdriverout 223.4e-3
rk1894 n1128__chipdriverout n1113__chipdriverout 142.4e-3
rk1895 n1113__chipdriverout n1114__chipdriverout 343.1e-3
rk1896 n1114__chipdriverout n1129__chipdriverout 239.6e-3
rk1897 n1129__chipdriverout n1117__chipdriverout 126.2e-3
rk1899 n1125__chipdriverout n1126__chipdriverout 3.1
rk1900 n1125__chipdriverout n1127__chipdriverout 3.1
rk1901 n1125__chipdriverout n1128__chipdriverout 3.1
rk1902 n1125__chipdriverout n1129__chipdriverout 3.1
rk1903 n15__i5__i7__xor2 n16__i5__i7__xor2 34.8e-3
rk1904 n2__i5__i7__xor2 n16__i5__i7__xor2 45
rk1905 n15__i5__i7__xor1 n16__i5__i7__xor1 34.8e-3
rk1906 n2__i5__i7__xor1 n16__i5__i7__xor1 45
rk1907 n394__i1__i14__net1 n509__i1__i14__net1 125e-3
rk1908 n396__i1__i14__net1 n510__i1__i14__net1 125e-3
rk1910 n650__vddio n652__vddio 30.13e-3
rk1911 n652__vddio n653__vddio 335.6e-3
rk1912 n653__vddio n654__vddio 343.1e-3
rk1913 n654__vddio n655__vddio 42.68e-3
rk1914 n655__vddio n656__vddio 321.2e-3
rk1915 n656__vddio n657__vddio 362.5e-3
rk1916 n657__vddio n658__vddio 40.17e-3
rk1917 n658__vddio n659__vddio 323.7e-3
rk1918 n659__vddio n660__vddio 343.1e-3
rk1919 n660__vddio n661__vddio 52.73e-3
rk1920 n661__vddio n662__vddio 394.2e-3
rk1921 n651__vddio n652__vddio 3.1
rk1922 n651__vddio n655__vddio 3.1
rk1923 n651__vddio n658__vddio 3.1
rk1924 n651__vddio n661__vddio 3.1
rk1925 n374__vss n371__vss 55.24e-3
rk1926 n371__vss n370__vss 365.7e-3
rk1927 n370__vss n375__vss 298.6e-3
rk1928 n375__vss n367__vss 42.68e-3
rk1929 n367__vss n366__vss 365.7e-3
rk1930 n366__vss n376__vss 187.7e-3
rk1931 n376__vss n377__vss 264.6e-3
rk1932 n373__vss n374__vss 3.75
rk1933 n373__vss n375__vss 3.75
rk1934 n373__vss n376__vss 5.7692
rk1935 n405__i1__i14__net1 n517__i1__i14__net1 125e-3
rk1936 n407__i1__i14__net1 n518__i1__i14__net1 125e-3
rk1938 n1133__chipdriverout n1134__chipdriverout 12.55e-3
rk1939 n1134__chipdriverout n1135__chipdriverout 365.7e-3
rk1940 n1135__chipdriverout n1136__chipdriverout 226.6e-3
rk1941 n1136__chipdriverout n1137__chipdriverout 116.5e-3
rk1942 n1137__chipdriverout n1138__chipdriverout 365.7e-3
rk1943 n1138__chipdriverout n1139__chipdriverout 242.8e-3
rk1944 n1139__chipdriverout n1140__chipdriverout 119.7e-3
rk1946 n1132__chipdriverout n1133__chipdriverout 5.7692
rk1947 n1132__chipdriverout n1136__chipdriverout 3.75
rk1948 n1132__chipdriverout n1139__chipdriverout 3.75
rk1950 n1143__chipdriverout n1145__chipdriverout 210.4e-3
rk1951 n1145__chipdriverout n1146__chipdriverout 155.3e-3
rk1952 n1146__chipdriverout n1147__chipdriverout 343.1e-3
rk1953 n1147__chipdriverout n1148__chipdriverout 226.6e-3
rk1954 n1148__chipdriverout n1149__chipdriverout 139.1e-3
rk1955 n1149__chipdriverout n1150__chipdriverout 362.5e-3
rk1956 n1150__chipdriverout n1151__chipdriverout 223.4e-3
rk1957 n1151__chipdriverout n1152__chipdriverout 142.4e-3
rk1958 n1152__chipdriverout n1153__chipdriverout 343.1e-3
rk1959 n1153__chipdriverout n1154__chipdriverout 239.6e-3
rk1960 n1154__chipdriverout n1155__chipdriverout 126.2e-3
rk1962 n1144__chipdriverout n1145__chipdriverout 3.1
rk1963 n1144__chipdriverout n1148__chipdriverout 3.1
rk1964 n1144__chipdriverout n1151__chipdriverout 3.1
rk1965 n1144__chipdriverout n1154__chipdriverout 3.1
rk1969 n671__vddio n686__vddio 30.13e-3
rk1970 n686__vddio n672__vddio 335.6e-3
rk1971 n672__vddio n675__vddio 343.1e-3
rk1972 n675__vddio n687__vddio 42.68e-3
rk1973 n687__vddio n676__vddio 321.2e-3
rk1974 n676__vddio n679__vddio 362.5e-3
rk1975 n679__vddio n688__vddio 40.17e-3
rk1976 n688__vddio n680__vddio 323.7e-3
rk1977 n680__vddio n683__vddio 343.1e-3
rk1978 n683__vddio n689__vddio 52.73e-3
rk1979 n689__vddio n690__vddio 394.2e-3
rk1980 n685__vddio n686__vddio 3.1
rk1981 n685__vddio n687__vddio 3.1
rk1982 n685__vddio n688__vddio 3.1
rk1983 n685__vddio n689__vddio 3.1
rk1984 n387__vss n384__vss 55.24e-3
rk1985 n384__vss n383__vss 365.7e-3
rk1986 n383__vss n388__vss 298.6e-3
rk1987 n388__vss n380__vss 42.68e-3
rk1988 n380__vss n379__vss 365.7e-3
rk1989 n379__vss n389__vss 187.7e-3
rk1990 n389__vss n390__vss 264.6e-3
rk1991 n386__vss n387__vss 3.75
rk1992 n386__vss n388__vss 3.75
rk1993 n386__vss n389__vss 5.7692
rk1994 n9__i5__i7__xor3 n11__i5__i7__xor3 10.91e-3
rk1995 n10__i5__i7__xor3 n11__i5__i7__xor3 31
rk1996 n9__i5__i7__xor0 n11__i5__i7__xor0 10.91e-3
rk1997 n10__i5__i7__xor0 n11__i5__i7__xor0 31
rk1998 n7__i5__i7__i5__net1 n8__i5__i7__i5__net1 31.2625
rk1999 n8__i5__i7__i5__net1 n9__i5__i7__i5__net1 75.1118
rk2000 n8__i5__i7__i5__net1 n3__i5__i7__i5__net1 213.9e-3
rk2001 n3__i5__i7__i5__net1 n10__i5__i7__i5__net1 125e-3
rk2002 n7__i5__i7__i4__net1 n8__i5__i7__i4__net1 31.2625
rk2003 n8__i5__i7__i4__net1 n9__i5__i7__i4__net1 75.1118
rk2004 n8__i5__i7__i4__net1 n3__i5__i7__i4__net1 213.9e-3
rk2005 n3__i5__i7__i4__net1 n10__i5__i7__i4__net1 125e-3
rk2006 n421__i1__i14__net1 n533__i1__i14__net1 125e-3
rk2007 n423__i1__i14__net1 n534__i1__i14__net1 125e-3
rk2009 n1172__chipdriverout n1173__chipdriverout 12.55e-3
rk2010 n1173__chipdriverout n1174__chipdriverout 365.7e-3
rk2011 n1174__chipdriverout n1175__chipdriverout 226.6e-3
rk2012 n1175__chipdriverout n1176__chipdriverout 116.5e-3
rk2013 n1176__chipdriverout n1177__chipdriverout 365.7e-3
rk2014 n1177__chipdriverout n1178__chipdriverout 242.8e-3
rk2015 n1178__chipdriverout n1179__chipdriverout 119.7e-3
rk2017 n1171__chipdriverout n1172__chipdriverout 5.7692
rk2018 n1171__chipdriverout n1175__chipdriverout 3.75
rk2019 n1171__chipdriverout n1178__chipdriverout 3.75
rk2021 n1182__chipdriverout n1184__chipdriverout 211.2e-3
rk2022 n1184__chipdriverout n1185__chipdriverout 156.2e-3
rk2023 n1185__chipdriverout n1186__chipdriverout 344.7e-3
rk2024 n1186__chipdriverout n1187__chipdriverout 227.4e-3
rk2025 n1187__chipdriverout n1188__chipdriverout 140e-3
rk2026 n1188__chipdriverout n1189__chipdriverout 364.2e-3
rk2027 n1189__chipdriverout n1190__chipdriverout 224.2e-3
rk2028 n1190__chipdriverout n1191__chipdriverout 143.2e-3
rk2029 n1191__chipdriverout n1192__chipdriverout 344.7e-3
rk2030 n1192__chipdriverout n1193__chipdriverout 240.4e-3
rk2031 n1193__chipdriverout n1194__chipdriverout 127e-3
rk2033 n1183__chipdriverout n1184__chipdriverout 3.1
rk2034 n1183__chipdriverout n1187__chipdriverout 3.1
rk2035 n1183__chipdriverout n1190__chipdriverout 3.1
rk2036 n1183__chipdriverout n1193__chipdriverout 3.1
rk2037 n8__i5__i7__net47 n7__i5__i7__net47 31.1227
rk2038 n7__i5__i7__net47 n9__i5__i7__net47 37.6081
rk2039 n6__i5__i7__net44 n4__i5__i7__net44 31.1227
rk2040 n4__i5__i7__net44 n7__i5__i7__net44 37.6081
rk2041 n426__i1__i14__net1 n537__i1__i14__net1 125e-3
rk2042 n428__i1__i14__net1 n538__i1__i14__net1 125e-3
rk2043 n392__vss n393__vss 55.24e-3
rk2044 n393__vss n394__vss 365.7e-3
rk2045 n394__vss n395__vss 298.6e-3
rk2046 n395__vss n396__vss 42.68e-3
rk2047 n396__vss n397__vss 365.7e-3
rk2048 n397__vss n398__vss 187.7e-3
rk2049 n398__vss n399__vss 264.6e-3
rk2050 n391__vss n392__vss 3.75
rk2051 n391__vss n395__vss 3.75
rk2052 n391__vss n398__vss 5.7692
rk2054 n692__vddio n694__vddio 30.13e-3
rk2055 n694__vddio n695__vddio 335.6e-3
rk2056 n695__vddio n696__vddio 343.1e-3
rk2057 n696__vddio n697__vddio 42.68e-3
rk2058 n697__vddio n698__vddio 321.2e-3
rk2059 n698__vddio n699__vddio 362.5e-3
rk2060 n699__vddio n700__vddio 40.17e-3
rk2061 n700__vddio n701__vddio 323.7e-3
rk2062 n701__vddio n702__vddio 343.1e-3
rk2063 n702__vddio n703__vddio 52.73e-3
rk2064 n703__vddio n704__vddio 394.2e-3
rk2065 n693__vddio n694__vddio 3.1
rk2066 n693__vddio n697__vddio 3.1
rk2067 n693__vddio n700__vddio 3.1
rk2068 n693__vddio n703__vddio 3.1
rk2069 n434__i1__i14__net1 n549__i1__i14__net1 125e-3
rk2070 n436__i1__i14__net1 n550__i1__i14__net1 125e-3
rk2071 n13__i5__i7__xor3 n14__i5__i7__xor3 4.428e-3
rk2072 n15__i5__i7__xor3 n16__i5__i7__xor3 4.428e-3
rk2073 n14__i5__i7__xor3 n16__i5__i7__xor3 15.28e-3
rk2074 n12__i5__i7__xor3 n13__i5__i7__xor3 75
rk2075 n13__i5__i7__xor0 n14__i5__i7__xor0 4.428e-3
rk2076 n15__i5__i7__xor0 n16__i5__i7__xor0 4.428e-3
rk2077 n14__i5__i7__xor0 n16__i5__i7__xor0 15.28e-3
rk2078 n12__i5__i7__xor0 n13__i5__i7__xor0 75
rk2080 n1211__chipdriverout n1212__chipdriverout 12.55e-3
rk2081 n1212__chipdriverout n1213__chipdriverout 365.7e-3
rk2082 n1213__chipdriverout n1214__chipdriverout 226.6e-3
rk2083 n1214__chipdriverout n1215__chipdriverout 116.5e-3
rk2084 n1215__chipdriverout n1216__chipdriverout 365.7e-3
rk2085 n1216__chipdriverout n1217__chipdriverout 242.8e-3
rk2086 n1217__chipdriverout n1218__chipdriverout 119.7e-3
rk2088 n1210__chipdriverout n1211__chipdriverout 5.7692
rk2089 n1210__chipdriverout n1214__chipdriverout 3.75
rk2090 n1210__chipdriverout n1217__chipdriverout 3.75
rk2092 n1221__chipdriverout n1223__chipdriverout 212.2e-3
rk2093 n1223__chipdriverout n1224__chipdriverout 157.2e-3
rk2094 n1224__chipdriverout n1225__chipdriverout 346.7e-3
rk2095 n1225__chipdriverout n1226__chipdriverout 228.4e-3
rk2096 n1226__chipdriverout n1227__chipdriverout 141e-3
rk2097 n1227__chipdriverout n1228__chipdriverout 366.1e-3
rk2098 n1228__chipdriverout n1229__chipdriverout 225.2e-3
rk2099 n1229__chipdriverout n1230__chipdriverout 144.2e-3
rk2100 n1230__chipdriverout n1231__chipdriverout 346.7e-3
rk2101 n1231__chipdriverout n1232__chipdriverout 241.4e-3
rk2102 n1232__chipdriverout n1233__chipdriverout 128e-3
rk2104 n1222__chipdriverout n1223__chipdriverout 3.1
rk2105 n1222__chipdriverout n1226__chipdriverout 3.1
rk2106 n1222__chipdriverout n1229__chipdriverout 3.1
rk2107 n1222__chipdriverout n1232__chipdriverout 3.1
rk2108 n442__i1__i14__net1 n557__i1__i14__net1 125e-3
rk2109 n444__i1__i14__net1 n558__i1__i14__net1 125e-3
rk2110 n405__vss n406__vss 55.24e-3
rk2111 n406__vss n407__vss 365.7e-3
rk2112 n407__vss n408__vss 298.6e-3
rk2113 n408__vss n409__vss 42.68e-3
rk2114 n409__vss n410__vss 365.7e-3
rk2115 n410__vss n411__vss 187.7e-3
rk2116 n411__vss n412__vss 264.6e-3
rk2117 n404__vss n405__vss 3.75
rk2118 n404__vss n408__vss 3.75
rk2119 n404__vss n411__vss 5.7692
rk2121 n713__vddio n715__vddio 30.13e-3
rk2122 n715__vddio n716__vddio 335.6e-3
rk2123 n716__vddio n717__vddio 343.1e-3
rk2124 n717__vddio n718__vddio 42.68e-3
rk2125 n718__vddio n719__vddio 321.2e-3
rk2126 n719__vddio n720__vddio 362.5e-3
rk2127 n720__vddio n721__vddio 40.17e-3
rk2128 n721__vddio n722__vddio 323.7e-3
rk2129 n722__vddio n723__vddio 343.1e-3
rk2130 n723__vddio n724__vddio 52.73e-3
rk2131 n724__vddio n725__vddio 394.2e-3
rk2132 n714__vddio n715__vddio 3.1
rk2133 n714__vddio n718__vddio 3.1
rk2134 n714__vddio n721__vddio 3.1
rk2135 n714__vddio n724__vddio 3.1
rk2136 n450__i1__i14__net1 n565__i1__i14__net1 125e-3
rk2137 n452__i1__i14__net1 n566__i1__i14__net1 125e-3
rk2139 n1250__chipdriverout n1251__chipdriverout 12.55e-3
rk2140 n1251__chipdriverout n1252__chipdriverout 365.7e-3
rk2141 n1252__chipdriverout n1253__chipdriverout 226.6e-3
rk2142 n1253__chipdriverout n1254__chipdriverout 116.5e-3
rk2143 n1254__chipdriverout n1255__chipdriverout 365.7e-3
rk2144 n1255__chipdriverout n1256__chipdriverout 242.8e-3
rk2145 n1256__chipdriverout n1257__chipdriverout 119.7e-3
rk2147 n1249__chipdriverout n1250__chipdriverout 5.7692
rk2148 n1249__chipdriverout n1253__chipdriverout 3.75
rk2149 n1249__chipdriverout n1256__chipdriverout 3.75
rk2151 n1260__chipdriverout n1262__chipdriverout 210.4e-3
rk2152 n1262__chipdriverout n1263__chipdriverout 155.3e-3
rk2153 n1263__chipdriverout n1264__chipdriverout 343.1e-3
rk2154 n1264__chipdriverout n1265__chipdriverout 226.6e-3
rk2155 n1265__chipdriverout n1266__chipdriverout 139.1e-3
rk2156 n1266__chipdriverout n1267__chipdriverout 362.5e-3
rk2157 n1267__chipdriverout n1268__chipdriverout 223.4e-3
rk2158 n1268__chipdriverout n1269__chipdriverout 142.4e-3
rk2159 n1269__chipdriverout n1270__chipdriverout 343.1e-3
rk2160 n1270__chipdriverout n1271__chipdriverout 239.6e-3
rk2161 n1271__chipdriverout n1272__chipdriverout 126.2e-3
rk2163 n1261__chipdriverout n1262__chipdriverout 3.1
rk2164 n1261__chipdriverout n1265__chipdriverout 3.1
rk2165 n1261__chipdriverout n1268__chipdriverout 3.1
rk2166 n1261__chipdriverout n1271__chipdriverout 3.1
rk2167 n9__i5__i7__net51 n10__i5__i7__net51 33.29e-3
rk2168 n10__i5__i7__net51 n8__i5__i7__net51 31.0291
rk2169 n8__i5__i7__net51 n9__i5__i7__net51 31
rk2170 n11__i5__i7__net51 n12__i5__i7__net51 75.0296
rk2171 n12__i5__i7__net51 n11__i5__i7__net51 75.0338
rk2172 n5__i5__i7__net50 n6__i5__i7__net50 33.29e-3
rk2173 n6__i5__i7__net50 n4__i5__i7__net50 31.0291
rk2174 n4__i5__i7__net50 n5__i5__i7__net50 31
rk2175 n7__i5__i7__net50 n8__i5__i7__net50 75.0296
rk2176 n8__i5__i7__net50 n7__i5__i7__net50 75.0338
rk2177 n458__i1__i14__net1 n573__i1__i14__net1 125e-3
rk2178 n460__i1__i14__net1 n574__i1__i14__net1 125e-3
rk2179 n14__i5__i7__xor2 n21__i5__i7__xor2 303.8e-3
rk2180 n21__i5__i7__xor2 n18__i5__i7__xor2 184.9e-3
rk2181 n18__i5__i7__xor2 n11__i5__i7__xor2 210.3e-3
rk2182 n21__i5__i7__xor2 n22__i5__i7__xor2 31.0934
rk2183 n14__i5__i7__xor1 n21__i5__i7__xor1 303.8e-3
rk2184 n21__i5__i7__xor1 n19__i5__i7__xor1 184.9e-3
rk2185 n19__i5__i7__xor1 n11__i5__i7__xor1 210.3e-3
rk2186 n21__i5__i7__xor1 n22__i5__i7__xor1 31.0934
rk2187 n6__i5__i7__i5__net1 n12__i5__i7__i5__net1 3.563e-3
rk2188 n12__i5__i7__i5__net1 n13__i5__i7__i5__net1 75.3952
rk2189 n6__i5__i7__i4__net1 n12__i5__i7__i4__net1 3.563e-3
rk2190 n12__i5__i7__i4__net1 n13__i5__i7__i4__net1 75.3952
rk2192 n734__vddio n736__vddio 30.13e-3
rk2193 n736__vddio n737__vddio 335.6e-3
rk2194 n737__vddio n738__vddio 343.1e-3
rk2195 n738__vddio n739__vddio 42.68e-3
rk2196 n739__vddio n740__vddio 321.2e-3
rk2197 n740__vddio n741__vddio 362.5e-3
rk2198 n741__vddio n742__vddio 40.17e-3
rk2199 n742__vddio n743__vddio 323.7e-3
rk2200 n743__vddio n744__vddio 343.1e-3
rk2201 n744__vddio n745__vddio 52.73e-3
rk2202 n745__vddio n746__vddio 394.2e-3
rk2203 n735__vddio n736__vddio 3.1
rk2204 n735__vddio n739__vddio 3.1
rk2205 n735__vddio n742__vddio 3.1
rk2206 n735__vddio n745__vddio 3.1
rk2207 n418__vss n419__vss 55.24e-3
rk2208 n419__vss n420__vss 365.7e-3
rk2209 n420__vss n421__vss 298.6e-3
rk2210 n421__vss n422__vss 42.68e-3
rk2211 n422__vss n423__vss 365.7e-3
rk2212 n423__vss n424__vss 187.7e-3
rk2213 n424__vss n425__vss 264.6e-3
rk2214 n417__vss n418__vss 3.75
rk2215 n417__vss n421__vss 3.75
rk2216 n417__vss n424__vss 5.7692
rk2217 n23__i5__i7__xor3 n24__i5__i7__xor3 31.115
rk2218 n24__i5__i7__xor3 n25__i5__i7__xor3 326.1e-3
rk2219 n25__i5__i7__xor3 n17__i5__i7__xor3 13.09e-3
rk2220 n24__i5__i7__xor3 n26__i5__i7__xor3 75.115
rk2221 n2__i5__i7__xor3 n25__i5__i7__xor3 15
rk2222 n23__i5__i7__xor0 n24__i5__i7__xor0 31.115
rk2223 n24__i5__i7__xor0 n25__i5__i7__xor0 326.1e-3
rk2224 n25__i5__i7__xor0 n17__i5__i7__xor0 13.09e-3
rk2225 n24__i5__i7__xor0 n26__i5__i7__xor0 75.115
rk2226 n2__i5__i7__xor0 n25__i5__i7__xor0 15
rk2227 n466__i1__i14__net1 n581__i1__i14__net1 125e-3
rk2228 n468__i1__i14__net1 n582__i1__i14__net1 125e-3
rk2230 n1289__chipdriverout n1290__chipdriverout 12.55e-3
rk2231 n1290__chipdriverout n1291__chipdriverout 365.7e-3
rk2232 n1291__chipdriverout n1292__chipdriverout 226.6e-3
rk2233 n1292__chipdriverout n1293__chipdriverout 116.5e-3
rk2234 n1293__chipdriverout n1294__chipdriverout 365.7e-3
rk2235 n1294__chipdriverout n1295__chipdriverout 242.8e-3
rk2236 n1295__chipdriverout n1296__chipdriverout 119.7e-3
rk2238 n1288__chipdriverout n1289__chipdriverout 5.7692
rk2239 n1288__chipdriverout n1292__chipdriverout 3.75
rk2240 n1288__chipdriverout n1295__chipdriverout 3.75
rk2242 n1299__chipdriverout n1301__chipdriverout 210.4e-3
rk2243 n1301__chipdriverout n1302__chipdriverout 155.3e-3
rk2244 n1302__chipdriverout n1303__chipdriverout 343.1e-3
rk2245 n1303__chipdriverout n1304__chipdriverout 226.6e-3
rk2246 n1304__chipdriverout n1305__chipdriverout 139.1e-3
rk2247 n1305__chipdriverout n1306__chipdriverout 362.5e-3
rk2248 n1306__chipdriverout n1307__chipdriverout 223.4e-3
rk2249 n1307__chipdriverout n1308__chipdriverout 142.4e-3
rk2250 n1308__chipdriverout n1309__chipdriverout 343.1e-3
rk2251 n1309__chipdriverout n1310__chipdriverout 239.6e-3
rk2252 n1310__chipdriverout n1311__chipdriverout 126.2e-3
rk2254 n1300__chipdriverout n1301__chipdriverout 3.1
rk2255 n1300__chipdriverout n1304__chipdriverout 3.1
rk2256 n1300__chipdriverout n1307__chipdriverout 3.1
rk2257 n1300__chipdriverout n1310__chipdriverout 3.1
rk2261 n755__vddio n757__vddio 30.13e-3
rk2262 n757__vddio n758__vddio 335.6e-3
rk2263 n758__vddio n759__vddio 343.1e-3
rk2264 n759__vddio n760__vddio 42.68e-3
rk2265 n760__vddio n761__vddio 321.2e-3
rk2266 n761__vddio n762__vddio 362.5e-3
rk2267 n762__vddio n763__vddio 40.17e-3
rk2268 n763__vddio n764__vddio 323.7e-3
rk2269 n764__vddio n765__vddio 343.1e-3
rk2270 n765__vddio n766__vddio 52.73e-3
rk2271 n766__vddio n767__vddio 394.2e-3
rk2272 n756__vddio n757__vddio 3.1
rk2273 n756__vddio n760__vddio 3.1
rk2274 n756__vddio n763__vddio 3.1
rk2275 n756__vddio n766__vddio 3.1
rk2276 n439__vss n437__vss 55.24e-3
rk2277 n437__vss n434__vss 365.7e-3
rk2278 n434__vss n440__vss 298.6e-3
rk2279 n440__vss n433__vss 42.68e-3
rk2280 n433__vss n430__vss 365.7e-3
rk2281 n430__vss n441__vss 187.7e-3
rk2282 n441__vss n442__vss 264.6e-3
rk2283 n438__vss n439__vss 3.75
rk2284 n438__vss n440__vss 3.75
rk2285 n438__vss n441__vss 5.7692
rk2286 n482__i1__i14__net1 n597__i1__i14__net1 125e-3
rk2287 n484__i1__i14__net1 n598__i1__i14__net1 125e-3
rk2288 n15__i5__i7__net51 n16__i5__i7__net51 34.8e-3
rk2289 n2__i5__i7__net51 n16__i5__i7__net51 45
rk2290 n2__i5__i7__net47 n10__i5__i7__net47 45.2869
rk2292 n1328__chipdriverout n1329__chipdriverout 12.55e-3
rk2293 n1329__chipdriverout n1330__chipdriverout 365.7e-3
rk2294 n1330__chipdriverout n1331__chipdriverout 226.6e-3
rk2295 n1331__chipdriverout n1332__chipdriverout 116.5e-3
rk2296 n1332__chipdriverout n1333__chipdriverout 365.7e-3
rk2297 n1333__chipdriverout n1334__chipdriverout 242.8e-3
rk2298 n1334__chipdriverout n1335__chipdriverout 119.7e-3
rk2300 n1327__chipdriverout n1328__chipdriverout 5.7692
rk2301 n1327__chipdriverout n1331__chipdriverout 3.75
rk2302 n1327__chipdriverout n1334__chipdriverout 3.75
rk2304 n1338__chipdriverout n1340__chipdriverout 211.2e-3
rk2305 n1340__chipdriverout n1341__chipdriverout 156.2e-3
rk2306 n1341__chipdriverout n1342__chipdriverout 344.7e-3
rk2307 n1342__chipdriverout n1343__chipdriverout 227.4e-3
rk2308 n1343__chipdriverout n1344__chipdriverout 140e-3
rk2309 n1344__chipdriverout n1345__chipdriverout 364.2e-3
rk2310 n1345__chipdriverout n1346__chipdriverout 224.2e-3
rk2311 n1346__chipdriverout n1347__chipdriverout 143.2e-3
rk2312 n1347__chipdriverout n1348__chipdriverout 344.7e-3
rk2313 n1348__chipdriverout n1349__chipdriverout 240.4e-3
rk2314 n1349__chipdriverout n1350__chipdriverout 127e-3
rk2316 n1339__chipdriverout n1340__chipdriverout 3.1
rk2317 n1339__chipdriverout n1343__chipdriverout 3.1
rk2318 n1339__chipdriverout n1346__chipdriverout 3.1
rk2319 n1339__chipdriverout n1349__chipdriverout 3.1
rk2320 n494__i1__i14__net1 n601__i1__i14__net1 125e-3
rk2321 n496__i1__i14__net1 n602__i1__i14__net1 125e-3
rk2323 n776__vddio n778__vddio 30.13e-3
rk2324 n778__vddio n779__vddio 335.6e-3
rk2325 n779__vddio n780__vddio 343.1e-3
rk2326 n780__vddio n781__vddio 42.68e-3
rk2327 n781__vddio n782__vddio 321.2e-3
rk2328 n782__vddio n783__vddio 362.5e-3
rk2329 n783__vddio n784__vddio 40.17e-3
rk2330 n784__vddio n785__vddio 323.7e-3
rk2331 n785__vddio n786__vddio 343.1e-3
rk2332 n786__vddio n787__vddio 52.73e-3
rk2333 n787__vddio n788__vddio 394.2e-3
rk2334 n777__vddio n778__vddio 3.1
rk2335 n777__vddio n781__vddio 3.1
rk2336 n777__vddio n784__vddio 3.1
rk2337 n777__vddio n787__vddio 3.1
rk2338 n444__vss n445__vss 55.24e-3
rk2339 n445__vss n446__vss 365.7e-3
rk2340 n446__vss n447__vss 298.6e-3
rk2341 n447__vss n448__vss 42.68e-3
rk2342 n448__vss n449__vss 365.7e-3
rk2343 n449__vss n450__vss 187.7e-3
rk2344 n450__vss n451__vss 264.6e-3
rk2345 n443__vss n444__vss 3.75
rk2346 n443__vss n447__vss 3.75
rk2347 n443__vss n450__vss 5.7692
rk2348 n498__i1__i14__net1 n613__i1__i14__net1 125e-3
rk2349 n500__i1__i14__net1 n614__i1__i14__net1 125e-3
rk2351 n1367__chipdriverout n1368__chipdriverout 12.55e-3
rk2352 n1368__chipdriverout n1369__chipdriverout 365.7e-3
rk2353 n1369__chipdriverout n1370__chipdriverout 226.6e-3
rk2354 n1370__chipdriverout n1371__chipdriverout 116.5e-3
rk2355 n1371__chipdriverout n1372__chipdriverout 365.7e-3
rk2356 n1372__chipdriverout n1373__chipdriverout 242.8e-3
rk2357 n1373__chipdriverout n1374__chipdriverout 119.7e-3
rk2359 n1366__chipdriverout n1367__chipdriverout 5.7692
rk2360 n1366__chipdriverout n1370__chipdriverout 3.75
rk2361 n1366__chipdriverout n1373__chipdriverout 3.75
rk2363 n1377__chipdriverout n1379__chipdriverout 210.4e-3
rk2364 n1379__chipdriverout n1380__chipdriverout 155.3e-3
rk2365 n1380__chipdriverout n1381__chipdriverout 343.1e-3
rk2366 n1381__chipdriverout n1382__chipdriverout 226.6e-3
rk2367 n1382__chipdriverout n1383__chipdriverout 139.1e-3
rk2368 n1383__chipdriverout n1384__chipdriverout 362.5e-3
rk2369 n1384__chipdriverout n1385__chipdriverout 223.4e-3
rk2370 n1385__chipdriverout n1386__chipdriverout 142.4e-3
rk2371 n1386__chipdriverout n1387__chipdriverout 343.1e-3
rk2372 n1387__chipdriverout n1388__chipdriverout 239.6e-3
rk2373 n1388__chipdriverout n1389__chipdriverout 126.2e-3
rk2375 n1378__chipdriverout n1379__chipdriverout 3.1
rk2376 n1378__chipdriverout n1382__chipdriverout 3.1
rk2377 n1378__chipdriverout n1385__chipdriverout 3.1
rk2378 n1378__chipdriverout n1388__chipdriverout 3.1
rk2379 n506__i1__i14__net1 n621__i1__i14__net1 125e-3
rk2380 n508__i1__i14__net1 n622__i1__i14__net1 125e-3
rk2381 n9__i5__i7__net50 n11__i5__i7__net50 10.91e-3
rk2382 n10__i5__i7__net50 n11__i5__i7__net50 31
rk2383 n9__i5__i7__i6__net1 n10__i5__i7__i6__net1 31.2625
rk2384 n10__i5__i7__i6__net1 n11__i5__i7__i6__net1 75.1118
rk2385 n10__i5__i7__i6__net1 n3__i5__i7__i6__net1 213.9e-3
rk2388 n801__vddio n803__vddio 30.13e-3
rk2389 n803__vddio n804__vddio 335.6e-3
rk2390 n804__vddio n805__vddio 343.1e-3
rk2391 n805__vddio n806__vddio 42.68e-3
rk2392 n806__vddio n807__vddio 321.2e-3
rk2393 n807__vddio n808__vddio 362.5e-3
rk2394 n808__vddio n809__vddio 40.17e-3
rk2395 n809__vddio n810__vddio 323.7e-3
rk2396 n810__vddio n811__vddio 343.1e-3
rk2397 n811__vddio n812__vddio 52.73e-3
rk2398 n812__vddio n813__vddio 394.2e-3
rk2399 n802__vddio n803__vddio 3.1
rk2400 n802__vddio n806__vddio 3.1
rk2401 n802__vddio n809__vddio 3.1
rk2402 n802__vddio n812__vddio 3.1
rk2403 n457__vss n458__vss 55.24e-3
rk2404 n458__vss n459__vss 365.7e-3
rk2405 n459__vss n460__vss 298.6e-3
rk2406 n460__vss n461__vss 42.68e-3
rk2407 n461__vss n462__vss 365.7e-3
rk2408 n462__vss n463__vss 187.7e-3
rk2409 n463__vss n464__vss 264.6e-3
rk2410 n456__vss n457__vss 3.75
rk2411 n456__vss n460__vss 3.75
rk2412 n456__vss n463__vss 5.7692
rk2413 n10__i5__i7__i7__net1 n11__i5__i7__i7__net1 33.29e-3
rk2414 n11__i5__i7__i7__net1 n9__i5__i7__i7__net1 31.0291
rk2415 n9__i5__i7__i7__net1 n10__i5__i7__i7__net1 31
rk2416 n12__i5__i7__i7__net1 n13__i5__i7__i7__net1 75.0296
rk2417 n13__i5__i7__i7__net1 n12__i5__i7__i7__net1 75.0338
rk2418 n514__i1__i14__net1 n625__i1__i14__net1 125e-3
rk2419 n516__i1__i14__net1 n626__i1__i14__net1 125e-3
rk2420 n6__i5__i7__net46 n4__i5__i7__net46 31.1227
rk2421 n4__i5__i7__net46 n7__i5__i7__net46 37.6081
rk2422 n3__i5__i7__i7__i0__net1 n5__i5__i7__i7__i0__net1 31.3722
rk2423 n5__i5__i7__i7__i0__net1 n7__i5__i7__i7__i0__net1 204.7e-3
rk2424 n7__i5__i7__i7__i0__net1 n2__i5__i7__i7__i0__net1 399.2e-3
rk2425 n4__i5__i7__i7__i0__net1 n5__i5__i7__i7__i0__net1 75
rk2426 n6__i5__i7__i7__i0__net1 n7__i5__i7__i7__i0__net1 75
rk2428 n1406__chipdriverout n1407__chipdriverout 12.55e-3
rk2429 n1407__chipdriverout n1408__chipdriverout 365.7e-3
rk2430 n1408__chipdriverout n1409__chipdriverout 226.6e-3
rk2431 n1409__chipdriverout n1410__chipdriverout 116.5e-3
rk2432 n1410__chipdriverout n1411__chipdriverout 365.7e-3
rk2433 n1411__chipdriverout n1412__chipdriverout 242.8e-3
rk2434 n1412__chipdriverout n1413__chipdriverout 119.7e-3
rk2436 n1405__chipdriverout n1406__chipdriverout 5.7692
rk2437 n1405__chipdriverout n1409__chipdriverout 3.75
rk2438 n1405__chipdriverout n1412__chipdriverout 3.75
rk2440 n1416__chipdriverout n1418__chipdriverout 210.4e-3
rk2441 n1418__chipdriverout n1419__chipdriverout 155.3e-3
rk2442 n1419__chipdriverout n1420__chipdriverout 343.1e-3
rk2443 n1420__chipdriverout n1421__chipdriverout 226.6e-3
rk2444 n1421__chipdriverout n1422__chipdriverout 139.1e-3
rk2445 n1422__chipdriverout n1423__chipdriverout 362.5e-3
rk2446 n1423__chipdriverout n1424__chipdriverout 223.4e-3
rk2447 n1424__chipdriverout n1425__chipdriverout 142.4e-3
rk2448 n1425__chipdriverout n1426__chipdriverout 343.1e-3
rk2449 n1426__chipdriverout n1427__chipdriverout 239.6e-3
rk2450 n1427__chipdriverout n1428__chipdriverout 126.2e-3
rk2452 n1417__chipdriverout n1418__chipdriverout 3.1
rk2453 n1417__chipdriverout n1421__chipdriverout 3.1
rk2454 n1417__chipdriverout n1424__chipdriverout 3.1
rk2455 n1417__chipdriverout n1427__chipdriverout 3.1
rk2456 n5__i5__i7__net47 n12__i5__i7__net47 292e-3
rk2457 n12__i5__i7__net47 n13__i5__i7__net47 31.1232
rk2458 n526__i1__i14__net1 n633__i1__i14__net1 125e-3
rk2459 n528__i1__i14__net1 n634__i1__i14__net1 125e-3
rk2460 n12__i5__i7__net44 n14__i5__i7__net44 9.718e-3
rk2461 n14__i5__i7__net44 n15__i5__i7__net44 115e-3
rk2462 n15__i5__i7__net44 n16__i5__i7__net44 328.8e-3
rk2463 n16__i5__i7__net44 n9__i5__i7__net44 11.8e-3
rk2464 n15__i5__i7__net44 n17__i5__i7__net44 75.115
rk2465 n13__i5__i7__net44 n14__i5__i7__net44 31
rk2466 n2__i5__i7__net44 n16__i5__i7__net44 15
rk2467 n13__i5__i7__net50 n14__i5__i7__net50 4.428e-3
rk2468 n15__i5__i7__net50 n16__i5__i7__net50 4.428e-3
rk2469 n14__i5__i7__net50 n16__i5__i7__net50 15.28e-3
rk2470 n12__i5__i7__net50 n13__i5__i7__net50 75
rk2472 n828__vddio n843__vddio 30.13e-3
rk2473 n843__vddio n829__vddio 335.6e-3
rk2474 n829__vddio n832__vddio 343.1e-3
rk2475 n832__vddio n844__vddio 42.68e-3
rk2476 n844__vddio n833__vddio 321.2e-3
rk2477 n833__vddio n836__vddio 362.5e-3
rk2478 n836__vddio n845__vddio 40.17e-3
rk2479 n845__vddio n837__vddio 323.7e-3
rk2480 n837__vddio n840__vddio 343.1e-3
rk2481 n840__vddio n846__vddio 52.73e-3
rk2482 n846__vddio n847__vddio 394.2e-3
rk2483 n842__vddio n843__vddio 3.1
rk2484 n842__vddio n844__vddio 3.1
rk2485 n842__vddio n845__vddio 3.1
rk2486 n842__vddio n846__vddio 3.1
rk2487 n478__vss n475__vss 55.24e-3
rk2488 n475__vss n474__vss 365.7e-3
rk2489 n474__vss n479__vss 298.6e-3
rk2490 n479__vss n471__vss 42.68e-3
rk2491 n471__vss n470__vss 365.7e-3
rk2492 n470__vss n480__vss 187.7e-3
rk2493 n480__vss n481__vss 264.6e-3
rk2494 n477__vss n478__vss 3.75
rk2495 n477__vss n479__vss 3.75
rk2496 n477__vss n480__vss 5.7692
rk2500 n1473__chipdriverout n1446__chipdriverout 12.55e-3
rk2501 n1446__chipdriverout n1447__chipdriverout 365.7e-3
rk2502 n1447__chipdriverout n1474__chipdriverout 226.6e-3
rk2503 n1474__chipdriverout n1450__chipdriverout 116.5e-3
rk2504 n1450__chipdriverout n1451__chipdriverout 365.7e-3
rk2505 n1451__chipdriverout n1475__chipdriverout 242.8e-3
rk2506 n1475__chipdriverout n1454__chipdriverout 119.7e-3
rk2508 n1472__chipdriverout n1473__chipdriverout 5.7692
rk2509 n1472__chipdriverout n1474__chipdriverout 3.75
rk2510 n1472__chipdriverout n1475__chipdriverout 3.75
rk2512 n1455__chipdriverout n1479__chipdriverout 210.4e-3
rk2513 n1479__chipdriverout n1458__chipdriverout 155.3e-3
rk2514 n1458__chipdriverout n1459__chipdriverout 343.1e-3
rk2515 n1459__chipdriverout n1480__chipdriverout 226.6e-3
rk2516 n1480__chipdriverout n1462__chipdriverout 139.1e-3
rk2517 n1462__chipdriverout n1463__chipdriverout 362.5e-3
rk2518 n1463__chipdriverout n1481__chipdriverout 223.4e-3
rk2519 n1481__chipdriverout n1466__chipdriverout 142.4e-3
rk2520 n1466__chipdriverout n1467__chipdriverout 343.1e-3
rk2521 n1467__chipdriverout n1482__chipdriverout 239.6e-3
rk2522 n1482__chipdriverout n1470__chipdriverout 126.2e-3
rk2524 n1478__chipdriverout n1479__chipdriverout 3.1
rk2525 n1478__chipdriverout n1480__chipdriverout 3.1
rk2526 n1478__chipdriverout n1481__chipdriverout 3.1
rk2527 n1478__chipdriverout n1482__chipdriverout 3.1
rk2528 n542__i1__i14__net1 n653__i1__i14__net1 125e-3
rk2529 n544__i1__i14__net1 n654__i1__i14__net1 125e-3
rk2531 n849__vddio n851__vddio 30.13e-3
rk2532 n851__vddio n852__vddio 335.6e-3
rk2533 n852__vddio n853__vddio 343.1e-3
rk2534 n853__vddio n854__vddio 42.68e-3
rk2535 n854__vddio n855__vddio 321.2e-3
rk2536 n855__vddio n856__vddio 362.5e-3
rk2537 n856__vddio n857__vddio 40.17e-3
rk2538 n857__vddio n858__vddio 323.7e-3
rk2539 n858__vddio n859__vddio 343.1e-3
rk2540 n859__vddio n860__vddio 52.73e-3
rk2541 n860__vddio n861__vddio 394.2e-3
rk2542 n850__vddio n851__vddio 3.1
rk2543 n850__vddio n854__vddio 3.1
rk2544 n850__vddio n857__vddio 3.1
rk2545 n850__vddio n860__vddio 3.1
rk2546 n483__vss n484__vss 55.24e-3
rk2547 n484__vss n485__vss 365.7e-3
rk2548 n485__vss n486__vss 298.6e-3
rk2549 n486__vss n487__vss 42.68e-3
rk2550 n487__vss n488__vss 365.7e-3
rk2551 n488__vss n489__vss 187.7e-3
rk2552 n489__vss n490__vss 264.6e-3
rk2553 n482__vss n483__vss 3.75
rk2554 n482__vss n486__vss 3.75
rk2555 n482__vss n489__vss 5.7692
rk2556 n2__i5__i7__i7__net1 n16__i5__i7__i7__net1 45.2869
rk2557 n546__i1__i14__net1 n661__i1__i14__net1 125e-3
rk2558 n548__i1__i14__net1 n662__i1__i14__net1 125e-3
rk2559 n5__i5__r0 n6__i5__r0 33.29e-3
rk2560 n6__i5__r0 n4__i5__r0 31.0291
rk2561 n4__i5__r0 n5__i5__r0 31
rk2562 n7__i5__r0 n8__i5__r0 75.0296
rk2563 n8__i5__r0 n7__i5__r0 75.0338
rk2565 n1500__chipdriverout n1501__chipdriverout 12.55e-3
rk2566 n1501__chipdriverout n1502__chipdriverout 365.7e-3
rk2567 n1502__chipdriverout n1503__chipdriverout 226.6e-3
rk2568 n1503__chipdriverout n1504__chipdriverout 116.5e-3
rk2569 n1504__chipdriverout n1505__chipdriverout 365.7e-3
rk2570 n1505__chipdriverout n1506__chipdriverout 242.8e-3
rk2571 n1506__chipdriverout n1507__chipdriverout 119.7e-3
rk2573 n1499__chipdriverout n1500__chipdriverout 5.7692
rk2574 n1499__chipdriverout n1503__chipdriverout 3.75
rk2575 n1499__chipdriverout n1506__chipdriverout 3.75
rk2577 n1510__chipdriverout n1512__chipdriverout 210.4e-3
rk2578 n1512__chipdriverout n1513__chipdriverout 155.3e-3
rk2579 n1513__chipdriverout n1514__chipdriverout 343.1e-3
rk2580 n1514__chipdriverout n1515__chipdriverout 226.6e-3
rk2581 n1515__chipdriverout n1516__chipdriverout 139.1e-3
rk2582 n1516__chipdriverout n1517__chipdriverout 362.5e-3
rk2583 n1517__chipdriverout n1518__chipdriverout 223.4e-3
rk2584 n1518__chipdriverout n1519__chipdriverout 142.4e-3
rk2585 n1519__chipdriverout n1520__chipdriverout 343.1e-3
rk2586 n1520__chipdriverout n1521__chipdriverout 239.6e-3
rk2587 n1521__chipdriverout n1522__chipdriverout 126.2e-3
rk2589 n1511__chipdriverout n1512__chipdriverout 3.1
rk2590 n1511__chipdriverout n1515__chipdriverout 3.1
rk2591 n1511__chipdriverout n1518__chipdriverout 3.1
rk2592 n1511__chipdriverout n1521__chipdriverout 3.1
rk2593 n7__i5__i7__net51 n21__i5__i7__net51 303.8e-3
rk2594 n21__i5__i7__net51 n18__i5__i7__net51 184.9e-3
rk2595 n18__i5__i7__net51 n4__i5__i7__net51 210.3e-3
rk2596 n21__i5__i7__net51 n22__i5__i7__net51 31.0934
rk2597 n6__i5__i7__i6__net1 n12__i5__i7__i6__net1 3.563e-3
rk2598 n12__i5__i7__i6__net1 n13__i5__i7__i6__net1 75.3952
rk2601 n21__i5__i7__net50 n22__i5__i7__net50 31.115
rk2602 n22__i5__i7__net50 n23__i5__i7__net50 326.1e-3
rk2603 n23__i5__i7__net50 n17__i5__i7__net50 13.09e-3
rk2604 n22__i5__i7__net50 n24__i5__i7__net50 75.115
rk2605 n2__i5__i7__net50 n23__i5__i7__net50 15
rk2607 n870__vddio n885__vddio 30.13e-3
rk2608 n885__vddio n871__vddio 335.6e-3
rk2609 n871__vddio n874__vddio 343.1e-3
rk2610 n874__vddio n886__vddio 42.68e-3
rk2611 n886__vddio n875__vddio 321.2e-3
rk2612 n875__vddio n878__vddio 362.5e-3
rk2613 n878__vddio n887__vddio 40.17e-3
rk2614 n887__vddio n879__vddio 323.7e-3
rk2615 n879__vddio n882__vddio 343.1e-3
rk2616 n882__vddio n888__vddio 52.73e-3
rk2617 n888__vddio n889__vddio 394.2e-3
rk2618 n884__vddio n885__vddio 3.1
rk2619 n884__vddio n886__vddio 3.1
rk2620 n884__vddio n887__vddio 3.1
rk2621 n884__vddio n888__vddio 3.1
rk2622 n504__vss n501__vss 55.24e-3
rk2623 n501__vss n500__vss 365.7e-3
rk2624 n500__vss n505__vss 298.6e-3
rk2625 n505__vss n497__vss 42.68e-3
rk2626 n497__vss n496__vss 365.7e-3
rk2627 n496__vss n506__vss 187.7e-3
rk2628 n506__vss n507__vss 264.6e-3
rk2629 n503__vss n504__vss 3.75
rk2630 n503__vss n505__vss 3.75
rk2631 n503__vss n506__vss 5.7692
rk2635 n1540__chipdriverout n1541__chipdriverout 12.55e-3
rk2636 n1541__chipdriverout n1542__chipdriverout 365.7e-3
rk2637 n1542__chipdriverout n1543__chipdriverout 226.6e-3
rk2638 n1543__chipdriverout n1544__chipdriverout 116.5e-3
rk2639 n1544__chipdriverout n1545__chipdriverout 365.7e-3
rk2640 n1545__chipdriverout n1546__chipdriverout 242.8e-3
rk2641 n1546__chipdriverout n1547__chipdriverout 119.7e-3
rk2643 n1539__chipdriverout n1540__chipdriverout 5.7692
rk2644 n1539__chipdriverout n1543__chipdriverout 3.75
rk2645 n1539__chipdriverout n1546__chipdriverout 3.75
rk2647 n1550__chipdriverout n1552__chipdriverout 210.4e-3
rk2648 n1552__chipdriverout n1553__chipdriverout 155.3e-3
rk2649 n1553__chipdriverout n1554__chipdriverout 343.1e-3
rk2650 n1554__chipdriverout n1555__chipdriverout 226.6e-3
rk2651 n1555__chipdriverout n1556__chipdriverout 139.1e-3
rk2652 n1556__chipdriverout n1557__chipdriverout 362.5e-3
rk2653 n1557__chipdriverout n1558__chipdriverout 223.4e-3
rk2654 n1558__chipdriverout n1559__chipdriverout 142.4e-3
rk2655 n1559__chipdriverout n1560__chipdriverout 343.1e-3
rk2656 n1560__chipdriverout n1561__chipdriverout 239.6e-3
rk2657 n1561__chipdriverout n1562__chipdriverout 126.2e-3
rk2659 n1551__chipdriverout n1552__chipdriverout 3.1
rk2660 n1551__chipdriverout n1555__chipdriverout 3.1
rk2661 n1551__chipdriverout n1558__chipdriverout 3.1
rk2662 n1551__chipdriverout n1561__chipdriverout 3.1
rk2663 n4__i5__clk_buf n17__i5__clk_buf 22.5251
rk2666 n2__i5__r1 n3__i5__r1 33.29e-3
rk2667 n3__i5__r1 i5__r1 31.0291
rk2668 i5__r1 n2__i5__r1 31
rk2669 n4__i5__r1 n5__i5__r1 75.0296
rk2670 n5__i5__r1 n4__i5__r1 75.0338
rk2672 n891__vddio n893__vddio 30.13e-3
rk2673 n893__vddio n894__vddio 335.6e-3
rk2674 n894__vddio n895__vddio 343.1e-3
rk2675 n895__vddio n896__vddio 42.68e-3
rk2676 n896__vddio n897__vddio 321.2e-3
rk2677 n897__vddio n898__vddio 362.5e-3
rk2678 n898__vddio n899__vddio 40.17e-3
rk2679 n899__vddio n900__vddio 323.7e-3
rk2680 n900__vddio n901__vddio 343.1e-3
rk2681 n901__vddio n902__vddio 52.73e-3
rk2682 n902__vddio n903__vddio 394.2e-3
rk2683 n892__vddio n893__vddio 3.1
rk2684 n892__vddio n896__vddio 3.1
rk2685 n892__vddio n899__vddio 3.1
rk2686 n892__vddio n902__vddio 3.1
rk2687 n509__vss n510__vss 55.24e-3
rk2688 n510__vss n511__vss 365.7e-3
rk2689 n511__vss n512__vss 298.6e-3
rk2690 n512__vss n513__vss 42.68e-3
rk2691 n513__vss n514__vss 365.7e-3
rk2692 n514__vss n515__vss 187.7e-3
rk2693 n515__vss n516__vss 264.6e-3
rk2694 n508__vss n509__vss 3.75
rk2695 n508__vss n512__vss 3.75
rk2696 n508__vss n515__vss 5.7692
rk2697 n3__i5__i7__i7__i1__net1 n5__i5__i7__i7__i1__net1 31.3722
rk2698 n5__i5__i7__i7__i1__net1 n7__i5__i7__i7__i1__net1 204.7e-3
rk2699 n7__i5__i7__i7__i1__net1 n2__i5__i7__i7__i1__net1 399.2e-3
rk2700 n4__i5__i7__i7__i1__net1 n5__i5__i7__i7__i1__net1 75
rk2701 n6__i5__i7__i7__i1__net1 n7__i5__i7__i7__i1__net1 75
rk2702 n5__i5__i7__i7__net1 n19__i5__i7__i7__net1 292e-3
rk2703 n19__i5__i7__i7__net1 n20__i5__i7__i7__net1 31.1232
rk2704 n578__i1__i14__net1 n693__i1__i14__net1 125e-3
rk2705 n580__i1__i14__net1 n694__i1__i14__net1 125e-3
rk2706 n14__i5__i7__net46 n15__i5__i7__net46 31.115
rk2707 n15__i5__i7__net46 n16__i5__i7__net46 328.8e-3
rk2708 n16__i5__i7__net46 n13__i5__i7__net46 11.8e-3
rk2709 n15__i5__i7__net46 n17__i5__i7__net46 75.115
rk2710 n2__i5__i7__net46 n16__i5__i7__net46 15
rk2712 n1580__chipdriverout n1581__chipdriverout 12.55e-3
rk2713 n1581__chipdriverout n1582__chipdriverout 365.7e-3
rk2714 n1582__chipdriverout n1583__chipdriverout 226.6e-3
rk2715 n1583__chipdriverout n1584__chipdriverout 116.5e-3
rk2716 n1584__chipdriverout n1585__chipdriverout 365.7e-3
rk2717 n1585__chipdriverout n1586__chipdriverout 242.8e-3
rk2718 n1586__chipdriverout n1587__chipdriverout 119.7e-3
rk2720 n1579__chipdriverout n1580__chipdriverout 5.7692
rk2721 n1579__chipdriverout n1583__chipdriverout 3.75
rk2722 n1579__chipdriverout n1586__chipdriverout 3.75
rk2724 n1590__chipdriverout n1592__chipdriverout 210.4e-3
rk2725 n1592__chipdriverout n1593__chipdriverout 155.3e-3
rk2726 n1593__chipdriverout n1594__chipdriverout 343.1e-3
rk2727 n1594__chipdriverout n1595__chipdriverout 226.6e-3
rk2728 n1595__chipdriverout n1596__chipdriverout 139.1e-3
rk2729 n1596__chipdriverout n1597__chipdriverout 362.5e-3
rk2730 n1597__chipdriverout n1598__chipdriverout 223.4e-3
rk2731 n1598__chipdriverout n1599__chipdriverout 142.4e-3
rk2732 n1599__chipdriverout n1600__chipdriverout 343.1e-3
rk2733 n1600__chipdriverout n1601__chipdriverout 239.6e-3
rk2734 n1601__chipdriverout n1602__chipdriverout 126.2e-3
rk2736 n1591__chipdriverout n1592__chipdriverout 3.1
rk2737 n1591__chipdriverout n1595__chipdriverout 3.1
rk2738 n1591__chipdriverout n1598__chipdriverout 3.1
rk2739 n1591__chipdriverout n1601__chipdriverout 3.1
rk2740 n8__i5__i6__net31 n9__i5__i6__net31 31.2664
rk2741 n9__i5__i6__net31 n10__i5__i6__net31 289.5e-3
rk2742 n10__i5__i6__net31 n11__i5__i6__net31 75.2422
rk2743 n9__i5__i6__net31 n12__i5__i6__net31 34.67e-3
rk2744 n12__i5__i6__net31 n13__i5__i6__net31 75.0632
rk2745 n10__i5__i6__net31 n14__i5__i6__net31 31.3039
rk2749 n922__vddio n924__vddio 30.13e-3
rk2750 n924__vddio n925__vddio 335.6e-3
rk2751 n925__vddio n926__vddio 343.1e-3
rk2752 n926__vddio n927__vddio 42.68e-3
rk2753 n927__vddio n928__vddio 321.2e-3
rk2754 n928__vddio n929__vddio 362.5e-3
rk2755 n929__vddio n930__vddio 40.17e-3
rk2756 n930__vddio n931__vddio 323.7e-3
rk2757 n931__vddio n932__vddio 343.1e-3
rk2758 n932__vddio n933__vddio 52.73e-3
rk2759 n933__vddio n934__vddio 394.2e-3
rk2760 n923__vddio n924__vddio 3.1
rk2761 n923__vddio n927__vddio 3.1
rk2762 n923__vddio n930__vddio 3.1
rk2763 n923__vddio n933__vddio 3.1
rk2764 n522__vss n523__vss 55.24e-3
rk2765 n523__vss n524__vss 365.7e-3
rk2766 n524__vss n525__vss 298.6e-3
rk2767 n525__vss n526__vss 42.68e-3
rk2768 n526__vss n527__vss 365.7e-3
rk2769 n527__vss n528__vss 187.7e-3
rk2770 n528__vss n529__vss 264.6e-3
rk2771 n521__vss n522__vss 3.75
rk2772 n521__vss n525__vss 3.75
rk2773 n521__vss n528__vss 5.7692
rk2775 n9__shift n2__shift 45.0049
rk2776 n594__i1__i14__net1 n709__i1__i14__net1 125e-3
rk2777 n596__i1__i14__net1 n710__i1__i14__net1 125e-3
rk2779 n1618__chipdriverout n1620__chipdriverout 210.4e-3
rk2780 n1620__chipdriverout n1621__chipdriverout 155.3e-3
rk2781 n1621__chipdriverout n1622__chipdriverout 343.1e-3
rk2782 n1622__chipdriverout n1623__chipdriverout 226.6e-3
rk2783 n1623__chipdriverout n1624__chipdriverout 139.1e-3
rk2784 n1624__chipdriverout n1625__chipdriverout 362.5e-3
rk2785 n1625__chipdriverout n1626__chipdriverout 223.4e-3
rk2786 n1626__chipdriverout n1627__chipdriverout 142.4e-3
rk2787 n1627__chipdriverout n1628__chipdriverout 343.1e-3
rk2788 n1628__chipdriverout n1629__chipdriverout 239.6e-3
rk2789 n1629__chipdriverout n1630__chipdriverout 126.2e-3
rk2791 n1619__chipdriverout n1620__chipdriverout 3.1
rk2792 n1619__chipdriverout n1623__chipdriverout 3.1
rk2793 n1619__chipdriverout n1626__chipdriverout 3.1
rk2794 n1619__chipdriverout n1629__chipdriverout 3.1
rk2796 n1634__chipdriverout n1635__chipdriverout 12.55e-3
rk2797 n1635__chipdriverout n1636__chipdriverout 365.7e-3
rk2798 n1636__chipdriverout n1637__chipdriverout 226.6e-3
rk2799 n1637__chipdriverout n1638__chipdriverout 116.5e-3
rk2800 n1638__chipdriverout n1639__chipdriverout 365.7e-3
rk2801 n1639__chipdriverout n1640__chipdriverout 242.8e-3
rk2802 n1640__chipdriverout n1641__chipdriverout 119.7e-3
rk2804 n1633__chipdriverout n1634__chipdriverout 5.7692
rk2805 n1633__chipdriverout n1637__chipdriverout 3.75
rk2806 n1633__chipdriverout n1640__chipdriverout 3.75
rk2807 n21__i5__i7__i7__net1 n26__i5__i7__i7__net1 38.44e-3
rk2808 n7__i5__i7__i7__net1 n26__i5__i7__i7__net1 45
rk2809 n606__i1__i14__net1 n717__i1__i14__net1 125e-3
rk2810 n608__i1__i14__net1 n718__i1__i14__net1 125e-3
rk2811 n43__vdd n44__vdd 31.2217
rk2812 n44__vdd n45__vdd 75.2494
rk2814 n943__vddio n945__vddio 30.13e-3
rk2815 n945__vddio n946__vddio 335.6e-3
rk2816 n946__vddio n947__vddio 343.1e-3
rk2817 n947__vddio n948__vddio 42.68e-3
rk2818 n948__vddio n949__vddio 321.2e-3
rk2819 n949__vddio n950__vddio 362.5e-3
rk2820 n950__vddio n951__vddio 40.17e-3
rk2821 n951__vddio n952__vddio 323.7e-3
rk2822 n952__vddio n953__vddio 343.1e-3
rk2823 n953__vddio n954__vddio 52.73e-3
rk2824 n954__vddio n955__vddio 394.2e-3
rk2825 n944__vddio n945__vddio 3.1
rk2826 n944__vddio n948__vddio 3.1
rk2827 n944__vddio n951__vddio 3.1
rk2828 n944__vddio n954__vddio 3.1
rk2829 n535__vss n536__vss 55.24e-3
rk2830 n536__vss n537__vss 365.7e-3
rk2831 n537__vss n538__vss 298.6e-3
rk2832 n538__vss n539__vss 42.68e-3
rk2833 n539__vss n540__vss 365.7e-3
rk2834 n540__vss n541__vss 187.7e-3
rk2835 n541__vss n542__vss 264.6e-3
rk2836 n534__vss n535__vss 3.75
rk2837 n534__vss n538__vss 3.75
rk2838 n534__vss n541__vss 5.7692
rk2839 n610__i1__i14__net1 n721__i1__i14__net1 125e-3
rk2840 n612__i1__i14__net1 n722__i1__i14__net1 125e-3
rk2842 n1657__chipdriverout n1659__chipdriverout 210.4e-3
rk2843 n1659__chipdriverout n1660__chipdriverout 155.3e-3
rk2844 n1660__chipdriverout n1661__chipdriverout 343.1e-3
rk2845 n1661__chipdriverout n1662__chipdriverout 226.6e-3
rk2846 n1662__chipdriverout n1663__chipdriverout 139.1e-3
rk2847 n1663__chipdriverout n1664__chipdriverout 362.5e-3
rk2848 n1664__chipdriverout n1665__chipdriverout 223.4e-3
rk2849 n1665__chipdriverout n1666__chipdriverout 142.4e-3
rk2850 n1666__chipdriverout n1667__chipdriverout 343.1e-3
rk2851 n1667__chipdriverout n1668__chipdriverout 239.6e-3
rk2852 n1668__chipdriverout n1669__chipdriverout 126.2e-3
rk2854 n1658__chipdriverout n1659__chipdriverout 3.1
rk2855 n1658__chipdriverout n1662__chipdriverout 3.1
rk2856 n1658__chipdriverout n1665__chipdriverout 3.1
rk2857 n1658__chipdriverout n1668__chipdriverout 3.1
rk2859 n1673__chipdriverout n1674__chipdriverout 12.55e-3
rk2860 n1674__chipdriverout n1675__chipdriverout 365.7e-3
rk2861 n1675__chipdriverout n1676__chipdriverout 226.6e-3
rk2862 n1676__chipdriverout n1677__chipdriverout 116.5e-3
rk2863 n1677__chipdriverout n1678__chipdriverout 365.7e-3
rk2864 n1678__chipdriverout n1679__chipdriverout 242.8e-3
rk2865 n1679__chipdriverout n1680__chipdriverout 119.7e-3
rk2867 n1672__chipdriverout n1673__chipdriverout 5.7692
rk2868 n1672__chipdriverout n1676__chipdriverout 3.75
rk2869 n1672__chipdriverout n1679__chipdriverout 3.75
rk2870 n618__i1__i14__net1 n725__i1__i14__net1 125e-3
rk2871 n620__i1__i14__net1 n726__i1__i14__net1 125e-3
rk2872 n3__i5__r2 n4__i5__r2 31.2117
rk2873 n4__i5__r2 n5__i5__r2 75.2117
rk2874 n4__i5__i6__i6__net4 n6__i5__i6__i6__net4 1.2154
rk2875 n6__i5__i6__i6__net4 n8__i5__i6__i6__net4 451.2e-3
rk2876 n8__i5__i6__i6__net4 n2__i5__i6__i6__net4 497.3e-3
rk2877 n5__i5__i6__i6__net4 n6__i5__i6__i6__net4 75
rk2878 n7__i5__i6__i6__net4 n8__i5__i6__i6__net4 31
rk2879 n7__shift n15__shift 1.3224
rk2880 n15__shift n5__shift 5.102e-3
rk2882 n964__vddio n966__vddio 30.13e-3
rk2883 n966__vddio n967__vddio 335.6e-3
rk2884 n967__vddio n968__vddio 343.1e-3
rk2885 n968__vddio n969__vddio 42.68e-3
rk2886 n969__vddio n970__vddio 321.2e-3
rk2887 n970__vddio n971__vddio 362.5e-3
rk2888 n971__vddio n972__vddio 40.17e-3
rk2889 n972__vddio n973__vddio 323.7e-3
rk2890 n973__vddio n974__vddio 343.1e-3
rk2891 n974__vddio n975__vddio 52.73e-3
rk2892 n975__vddio n976__vddio 394.2e-3
rk2893 n965__vddio n966__vddio 3.1
rk2894 n965__vddio n969__vddio 3.1
rk2895 n965__vddio n972__vddio 3.1
rk2896 n965__vddio n975__vddio 3.1
rk2897 n554__vss n555__vss 55.24e-3
rk2898 n555__vss n556__vss 365.7e-3
rk2899 n556__vss n557__vss 298.6e-3
rk2900 n557__vss n558__vss 42.68e-3
rk2901 n558__vss n559__vss 365.7e-3
rk2902 n559__vss n560__vss 187.7e-3
rk2903 n560__vss n561__vss 264.6e-3
rk2904 n553__vss n554__vss 3.75
rk2905 n553__vss n557__vss 3.75
rk2906 n553__vss n560__vss 5.7692
rk2907 n8__i5__i6__net30 n9__i5__i6__net30 75.2457
rk2908 n9__i5__i6__net30 n11__i5__i6__net30 219e-3
rk2909 n11__i5__i6__net30 n13__i5__i6__net30 1.1197
rk2910 n13__i5__i6__net30 n14__i5__i6__net30 75.5378
rk2911 n10__i5__i6__net30 n11__i5__i6__net30 31
rk2912 n12__i5__i6__net30 n13__i5__i6__net30 31
rk2913 n11__i5__i7__net44 n21__i5__i7__net44 250e-3
rk2914 n630__i1__i14__net1 n729__i1__i14__net1 125e-3
rk2915 n632__i1__i14__net1 n730__i1__i14__net1 125e-3
rk2917 n1696__chipdriverout n1698__chipdriverout 210.4e-3
rk2918 n1698__chipdriverout n1699__chipdriverout 155.3e-3
rk2919 n1699__chipdriverout n1700__chipdriverout 343.1e-3
rk2920 n1700__chipdriverout n1701__chipdriverout 226.6e-3
rk2921 n1701__chipdriverout n1702__chipdriverout 139.1e-3
rk2922 n1702__chipdriverout n1703__chipdriverout 362.5e-3
rk2923 n1703__chipdriverout n1704__chipdriverout 223.4e-3
rk2924 n1704__chipdriverout n1705__chipdriverout 142.4e-3
rk2925 n1705__chipdriverout n1706__chipdriverout 343.1e-3
rk2926 n1706__chipdriverout n1707__chipdriverout 239.6e-3
rk2927 n1707__chipdriverout n1708__chipdriverout 126.2e-3
rk2929 n1697__chipdriverout n1698__chipdriverout 3.1
rk2930 n1697__chipdriverout n1701__chipdriverout 3.1
rk2931 n1697__chipdriverout n1704__chipdriverout 3.1
rk2932 n1697__chipdriverout n1707__chipdriverout 3.1
rk2934 n1712__chipdriverout n1713__chipdriverout 12.55e-3
rk2935 n1713__chipdriverout n1714__chipdriverout 365.7e-3
rk2936 n1714__chipdriverout n1715__chipdriverout 226.6e-3
rk2937 n1715__chipdriverout n1716__chipdriverout 116.5e-3
rk2938 n1716__chipdriverout n1717__chipdriverout 365.7e-3
rk2939 n1717__chipdriverout n1718__chipdriverout 242.8e-3
rk2940 n1718__chipdriverout n1719__chipdriverout 119.7e-3
rk2942 n1711__chipdriverout n1712__chipdriverout 5.7692
rk2943 n1711__chipdriverout n1715__chipdriverout 3.75
rk2944 n1711__chipdriverout n1718__chipdriverout 3.75
rk2945 n2__i5__i6__i2__net25 n3__i5__i6__i2__net25 323.3e-3
rk2946 i5__i6__i2__net25 n2__i5__i6__i2__net25 15.5
rk2947 i5__i6__i2__net21 n2__i5__i6__i2__net21 37.7516
rk2948 n638__i1__i14__net1 n733__i1__i14__net1 125e-3
rk2949 n640__i1__i14__net1 n734__i1__i14__net1 125e-3
rk2950 n5__i5__i7__i7__net2 n6__i5__i7__i7__net2 31.2168
rk2951 n6__i5__i7__i7__net2 n7__i5__i7__i7__net2 75.1565
rk2952 n6__i5__i7__i7__net2 n8__i5__i7__i7__net2 440.6e-3
rk2953 n8__i5__i7__i7__net2 n4__i5__i7__i7__net2 227.3e-3
rk2954 n8__i5__i7__i7__net2 n2__i5__i7__i7__net2 44.01e-3
rk2955 n9__i5__i7__net46 n18__i5__i7__net46 250e-3
rk2956 n3__i5__i6__net30 n15__i5__i6__net30 22.8737
rk2958 n985__vddio n987__vddio 30.13e-3
rk2959 n987__vddio n988__vddio 335.6e-3
rk2960 n988__vddio n989__vddio 343.1e-3
rk2961 n989__vddio n990__vddio 42.68e-3
rk2962 n990__vddio n991__vddio 321.2e-3
rk2963 n991__vddio n992__vddio 362.5e-3
rk2964 n992__vddio n993__vddio 40.17e-3
rk2965 n993__vddio n994__vddio 323.7e-3
rk2966 n994__vddio n995__vddio 343.1e-3
rk2967 n995__vddio n996__vddio 52.73e-3
rk2968 n996__vddio n997__vddio 394.2e-3
rk2969 n986__vddio n987__vddio 3.1
rk2970 n986__vddio n990__vddio 3.1
rk2971 n986__vddio n993__vddio 3.1
rk2972 n986__vddio n996__vddio 3.1
rk2973 n567__vss n568__vss 55.24e-3
rk2974 n568__vss n569__vss 365.7e-3
rk2975 n569__vss n570__vss 298.6e-3
rk2976 n570__vss n571__vss 42.68e-3
rk2977 n571__vss n572__vss 365.7e-3
rk2978 n572__vss n573__vss 187.7e-3
rk2979 n573__vss n574__vss 264.6e-3
rk2980 n566__vss n567__vss 3.75
rk2981 n566__vss n570__vss 3.75
rk2982 n566__vss n573__vss 5.7692
rk2983 n4__i5__i7__i7__net3 n6__i5__i7__i7__net3 31.0041
rk2985 n6__i5__i7__i7__net3 n4__i5__i7__i7__net3 31.0038
rk2986 n5__i5__i7__i7__net3 n6__i5__i7__i7__net3 37.5
rk2987 n5__i5__i6__i2__net25 n6__i5__i6__i2__net25 350.8e-3
rk2988 n4__i5__i6__i2__net25 n5__i5__i6__i2__net25 15.5
rk2989 n3__i5__i6__i2__net21 n5__i5__i6__i2__net21 4.9e-3
rk2990 n4__i5__i6__i2__net21 n5__i5__i6__i2__net21 37.5
rk2991 n646__i1__i14__net1 n737__i1__i14__net1 125e-3
rk2992 n648__i1__i14__net1 n738__i1__i14__net1 125e-3
rk2993 n3__i5__i6__net31 n17__i5__i6__net31 500e-3
rk2996 n1735__chipdriverout n1737__chipdriverout 210.4e-3
rk2997 n1737__chipdriverout n1738__chipdriverout 155.3e-3
rk2998 n1738__chipdriverout n1739__chipdriverout 343.1e-3
rk2999 n1739__chipdriverout n1740__chipdriverout 226.6e-3
rk3000 n1740__chipdriverout n1741__chipdriverout 139.1e-3
rk3001 n1741__chipdriverout n1742__chipdriverout 362.5e-3
rk3002 n1742__chipdriverout n1743__chipdriverout 223.4e-3
rk3003 n1743__chipdriverout n1744__chipdriverout 142.4e-3
rk3004 n1744__chipdriverout n1745__chipdriverout 343.1e-3
rk3005 n1745__chipdriverout n1746__chipdriverout 239.6e-3
rk3006 n1746__chipdriverout n1747__chipdriverout 126.2e-3
rk3008 n1736__chipdriverout n1737__chipdriverout 3.1
rk3009 n1736__chipdriverout n1740__chipdriverout 3.1
rk3010 n1736__chipdriverout n1743__chipdriverout 3.1
rk3011 n1736__chipdriverout n1746__chipdriverout 3.1
rk3013 n1751__chipdriverout n1752__chipdriverout 12.55e-3
rk3014 n1752__chipdriverout n1753__chipdriverout 365.7e-3
rk3015 n1753__chipdriverout n1754__chipdriverout 226.6e-3
rk3016 n1754__chipdriverout n1755__chipdriverout 116.5e-3
rk3017 n1755__chipdriverout n1756__chipdriverout 365.7e-3
rk3018 n1756__chipdriverout n1757__chipdriverout 242.8e-3
rk3019 n1757__chipdriverout n1758__chipdriverout 119.7e-3
rk3021 n1750__chipdriverout n1751__chipdriverout 5.7692
rk3022 n1750__chipdriverout n1754__chipdriverout 3.75
rk3023 n1750__chipdriverout n1757__chipdriverout 3.75
rk3024 n10__i5__i7__net46 n23__i5__i7__net46 250e-3
rk3025 n650__i1__i14__net1 n741__i1__i14__net1 125e-3
rk3026 n652__i1__i14__net1 n742__i1__i14__net1 125e-3
rk3027 n8__i5__i6__i2__net25 n9__i5__i6__i2__net25 350.8e-3
rk3028 n7__i5__i6__i2__net25 n8__i5__i6__i2__net25 15.5
rk3029 n6__i5__i6__i2__net21 n8__i5__i6__i2__net21 4.9e-3
rk3030 n7__i5__i6__i2__net21 n8__i5__i6__i2__net21 37.5
rk3032 n1005__vddio n1021__vddio 30.13e-3
rk3033 n1021__vddio n1008__vddio 335.6e-3
rk3034 n1008__vddio n1009__vddio 343.1e-3
rk3035 n1009__vddio n1022__vddio 42.68e-3
rk3036 n1022__vddio n1012__vddio 321.2e-3
rk3037 n1012__vddio n1013__vddio 362.5e-3
rk3038 n1013__vddio n1023__vddio 40.17e-3
rk3039 n1023__vddio n1016__vddio 323.7e-3
rk3040 n1016__vddio n1017__vddio 343.1e-3
rk3041 n1017__vddio n1024__vddio 52.73e-3
rk3042 n1024__vddio n1025__vddio 394.2e-3
rk3043 n1020__vddio n1021__vddio 3.1
rk3044 n1020__vddio n1022__vddio 3.1
rk3045 n1020__vddio n1023__vddio 3.1
rk3046 n1020__vddio n1024__vddio 3.1
rk3047 n588__vss n586__vss 55.24e-3
rk3048 n586__vss n583__vss 365.7e-3
rk3049 n583__vss n589__vss 298.6e-3
rk3050 n589__vss n582__vss 42.68e-3
rk3051 n582__vss n579__vss 365.7e-3
rk3052 n579__vss n590__vss 187.7e-3
rk3053 n590__vss n591__vss 264.6e-3
rk3054 n587__vss n588__vss 3.75
rk3055 n587__vss n589__vss 3.75
rk3056 n587__vss n590__vss 5.7692
rk3057 n14__i5__i7__i7__net1 n27__i5__i7__i7__net1 241.6e-3
rk3058 n27__i5__i7__i7__net1 n17__i5__i7__i7__net1 6.874e-3
rk3060 n658__i1__i14__net1 n745__i1__i14__net1 125e-3
rk3061 n660__i1__i14__net1 n746__i1__i14__net1 125e-3
rk3062 n2__i5__i6__i2__net24 n3__i5__i6__i2__net24 323.3e-3
rk3063 i5__i6__i2__net24 n2__i5__i6__i2__net24 15.5
rk3064 i5__i6__i2__net23 n2__i5__i6__i2__net23 37.7516
rk3066 n1774__chipdriverout n1776__chipdriverout 210.4e-3
rk3067 n1776__chipdriverout n1777__chipdriverout 155.3e-3
rk3068 n1777__chipdriverout n1778__chipdriverout 343.1e-3
rk3069 n1778__chipdriverout n1779__chipdriverout 226.6e-3
rk3070 n1779__chipdriverout n1780__chipdriverout 139.1e-3
rk3071 n1780__chipdriverout n1781__chipdriverout 362.5e-3
rk3072 n1781__chipdriverout n1782__chipdriverout 223.4e-3
rk3073 n1782__chipdriverout n1783__chipdriverout 142.4e-3
rk3074 n1783__chipdriverout n1784__chipdriverout 343.1e-3
rk3075 n1784__chipdriverout n1785__chipdriverout 239.6e-3
rk3076 n1785__chipdriverout n1786__chipdriverout 126.2e-3
rk3078 n1775__chipdriverout n1776__chipdriverout 3.1
rk3079 n1775__chipdriverout n1779__chipdriverout 3.1
rk3080 n1775__chipdriverout n1782__chipdriverout 3.1
rk3081 n1775__chipdriverout n1785__chipdriverout 3.1
rk3083 n1790__chipdriverout n1791__chipdriverout 12.55e-3
rk3084 n1791__chipdriverout n1792__chipdriverout 365.7e-3
rk3085 n1792__chipdriverout n1793__chipdriverout 226.6e-3
rk3086 n1793__chipdriverout n1794__chipdriverout 116.5e-3
rk3087 n1794__chipdriverout n1795__chipdriverout 365.7e-3
rk3088 n1795__chipdriverout n1796__chipdriverout 242.8e-3
rk3089 n1796__chipdriverout n1797__chipdriverout 119.7e-3
rk3091 n1789__chipdriverout n1790__chipdriverout 5.7692
rk3092 n1789__chipdriverout n1793__chipdriverout 3.75
rk3093 n1789__chipdriverout n1796__chipdriverout 3.75
rk3094 n8__i5__i6__i2__net22 n9__i5__i6__i2__net22 15.9814
rk3095 n9__i5__i6__i2__net22 n10__i5__i6__i2__net22 37.8249
rk3096 n9__i5__i6__i2__net22 n3__i5__i6__i2__net22 22.9156
rk3097 n670__i1__i14__net1 n749__i1__i14__net1 125e-3
rk3098 n672__i1__i14__net1 n750__i1__i14__net1 125e-3
rk3099 n5__i5__i6__i2__net24 n6__i5__i6__i2__net24 350.8e-3
rk3100 n4__i5__i6__i2__net24 n5__i5__i6__i2__net24 15.5
rk3101 n3__i5__i6__i2__net23 n5__i5__i6__i2__net23 4.9e-3
rk3102 n4__i5__i6__i2__net23 n5__i5__i6__i2__net23 37.5
rk3104 n1037__vddio n1039__vddio 30.13e-3
rk3105 n1039__vddio n1040__vddio 335.6e-3
rk3106 n1040__vddio n1041__vddio 343.1e-3
rk3107 n1041__vddio n1042__vddio 42.68e-3
rk3108 n1042__vddio n1043__vddio 321.2e-3
rk3109 n1043__vddio n1044__vddio 362.5e-3
rk3110 n1044__vddio n1045__vddio 40.17e-3
rk3111 n1045__vddio n1046__vddio 323.7e-3
rk3112 n1046__vddio n1047__vddio 343.1e-3
rk3113 n1047__vddio n1048__vddio 52.73e-3
rk3114 n1048__vddio n1049__vddio 394.2e-3
rk3115 n1038__vddio n1039__vddio 3.1
rk3116 n1038__vddio n1042__vddio 3.1
rk3117 n1038__vddio n1045__vddio 3.1
rk3118 n1038__vddio n1048__vddio 3.1
rk3119 n593__vss n594__vss 55.24e-3
rk3120 n594__vss n595__vss 365.7e-3
rk3121 n595__vss n596__vss 298.6e-3
rk3122 n596__vss n597__vss 42.68e-3
rk3123 n597__vss n598__vss 365.7e-3
rk3124 n598__vss n599__vss 187.7e-3
rk3125 n599__vss n600__vss 264.6e-3
rk3126 n592__vss n593__vss 3.75
rk3127 n592__vss n596__vss 3.75
rk3128 n592__vss n599__vss 5.7692
rk3130 n15__i5__clk_buf n35__i5__clk_buf 500e-3
rk3131 n2__i5__i7__i7__net3 n8__i5__i7__i7__net3 45.2925
rk3132 n674__i1__i14__net1 n753__i1__i14__net1 125e-3
rk3133 n676__i1__i14__net1 n754__i1__i14__net1 125e-3
rk3134 n8__i5__i6__i2__net24 n9__i5__i6__i2__net24 350.8e-3
rk3135 n7__i5__i6__i2__net24 n8__i5__i6__i2__net24 15.5
rk3136 n6__i5__i6__i2__net23 n8__i5__i6__i2__net23 4.9e-3
rk3137 n7__i5__i6__i2__net23 n8__i5__i6__i2__net23 37.5
rk3139 n1824__chipdriverout n1812__chipdriverout 12.55e-3
rk3140 n1812__chipdriverout n1815__chipdriverout 365.7e-3
rk3141 n1815__chipdriverout n1825__chipdriverout 226.6e-3
rk3142 n1825__chipdriverout n1816__chipdriverout 116.5e-3
rk3143 n1816__chipdriverout n1819__chipdriverout 365.7e-3
rk3144 n1819__chipdriverout n1826__chipdriverout 242.8e-3
rk3145 n1826__chipdriverout n1820__chipdriverout 119.7e-3
rk3147 n1823__chipdriverout n1824__chipdriverout 5.7692
rk3148 n1823__chipdriverout n1825__chipdriverout 3.75
rk3149 n1823__chipdriverout n1826__chipdriverout 3.75
rk3151 n1829__chipdriverout n1831__chipdriverout 210.4e-3
rk3152 n1831__chipdriverout n1832__chipdriverout 155.3e-3
rk3153 n1832__chipdriverout n1833__chipdriverout 343.1e-3
rk3154 n1833__chipdriverout n1834__chipdriverout 226.6e-3
rk3155 n1834__chipdriverout n1835__chipdriverout 139.1e-3
rk3156 n1835__chipdriverout n1836__chipdriverout 362.5e-3
rk3157 n1836__chipdriverout n1837__chipdriverout 223.4e-3
rk3158 n1837__chipdriverout n1838__chipdriverout 142.4e-3
rk3159 n1838__chipdriverout n1839__chipdriverout 343.1e-3
rk3160 n1839__chipdriverout n1840__chipdriverout 239.6e-3
rk3161 n1840__chipdriverout n1841__chipdriverout 126.2e-3
rk3163 n1830__chipdriverout n1831__chipdriverout 3.1
rk3164 n1830__chipdriverout n1834__chipdriverout 3.1
rk3165 n1830__chipdriverout n1837__chipdriverout 3.1
rk3166 n1830__chipdriverout n1840__chipdriverout 3.1
rk3167 n10__i5__r2 n9__i5__r2 31.1111
rk3168 n9__i5__r2 n11__i5__r2 75.2193
rk3171 n38__reset n40__reset 250e-3
rk3173 n1058__vddio n1060__vddio 30.13e-3
rk3174 n1060__vddio n1061__vddio 335.6e-3
rk3175 n1061__vddio n1062__vddio 343.1e-3
rk3176 n1062__vddio n1063__vddio 42.68e-3
rk3177 n1063__vddio n1064__vddio 321.2e-3
rk3178 n1064__vddio n1065__vddio 362.5e-3
rk3179 n1065__vddio n1066__vddio 40.17e-3
rk3180 n1066__vddio n1067__vddio 323.7e-3
rk3181 n1067__vddio n1068__vddio 343.1e-3
rk3182 n1068__vddio n1069__vddio 52.73e-3
rk3183 n1069__vddio n1070__vddio 394.2e-3
rk3184 n1059__vddio n1060__vddio 3.1
rk3185 n1059__vddio n1063__vddio 3.1
rk3186 n1059__vddio n1066__vddio 3.1
rk3187 n1059__vddio n1069__vddio 3.1
rk3188 n606__vss n607__vss 55.24e-3
rk3189 n607__vss n608__vss 365.7e-3
rk3190 n608__vss n609__vss 298.6e-3
rk3191 n609__vss n610__vss 42.68e-3
rk3192 n610__vss n611__vss 365.7e-3
rk3193 n611__vss n612__vss 187.7e-3
rk3194 n612__vss n613__vss 264.6e-3
rk3195 n605__vss n606__vss 3.75
rk3196 n605__vss n609__vss 3.75
rk3197 n605__vss n612__vss 5.7692
rk3200 n4__clk_out n8__clk_out 45.2798
rk3202 n1852__chipdriverout n1854__chipdriverout 210.4e-3
rk3203 n1854__chipdriverout n1855__chipdriverout 155.3e-3
rk3204 n1855__chipdriverout n1856__chipdriverout 343.1e-3
rk3205 n1856__chipdriverout n1857__chipdriverout 226.6e-3
rk3206 n1857__chipdriverout n1858__chipdriverout 139.1e-3
rk3207 n1858__chipdriverout n1859__chipdriverout 362.5e-3
rk3208 n1859__chipdriverout n1860__chipdriverout 223.4e-3
rk3209 n1860__chipdriverout n1861__chipdriverout 142.4e-3
rk3210 n1861__chipdriverout n1862__chipdriverout 343.1e-3
rk3211 n1862__chipdriverout n1863__chipdriverout 239.6e-3
rk3212 n1863__chipdriverout n1864__chipdriverout 126.2e-3
rk3214 n1853__chipdriverout n1854__chipdriverout 3.1
rk3215 n1853__chipdriverout n1857__chipdriverout 3.1
rk3216 n1853__chipdriverout n1860__chipdriverout 3.1
rk3217 n1853__chipdriverout n1863__chipdriverout 3.1
rk3219 n1868__chipdriverout n1869__chipdriverout 12.55e-3
rk3220 n1869__chipdriverout n1870__chipdriverout 365.7e-3
rk3221 n1870__chipdriverout n1871__chipdriverout 226.6e-3
rk3222 n1871__chipdriverout n1872__chipdriverout 116.5e-3
rk3223 n1872__chipdriverout n1873__chipdriverout 365.7e-3
rk3224 n1873__chipdriverout n1874__chipdriverout 242.8e-3
rk3225 n1874__chipdriverout n1875__chipdriverout 119.7e-3
rk3227 n1867__chipdriverout n1868__chipdriverout 5.7692
rk3228 n1867__chipdriverout n1871__chipdriverout 3.75
rk3229 n1867__chipdriverout n1874__chipdriverout 3.75
rk3230 i5__i6__net32 n2__i5__i6__net32 19.0609
rk3231 n2__i5__i6__net32 n3__i5__i6__net32 293e-3
rk3232 n3__i5__i6__net32 n4__i5__i6__net32 420.4e-3
rk3233 n4__i5__i6__net32 n5__i5__i6__net32 37.828
rk3234 n3__i5__i6__net32 n6__i5__i6__net32 19.0309
rk3235 n4__i5__i6__net32 n7__i5__i6__net32 15.8422
rk3236 n702__i1__i14__net1 n765__i1__i14__net1 125e-3
rk3237 n704__i1__i14__net1 n766__i1__i14__net1 125e-3
rk3239 n1079__vddio n1081__vddio 30.13e-3
rk3240 n1081__vddio n1082__vddio 335.6e-3
rk3241 n1082__vddio n1083__vddio 343.1e-3
rk3242 n1083__vddio n1084__vddio 42.68e-3
rk3243 n1084__vddio n1085__vddio 321.2e-3
rk3244 n1085__vddio n1086__vddio 362.5e-3
rk3245 n1086__vddio n1087__vddio 40.17e-3
rk3246 n1087__vddio n1088__vddio 323.7e-3
rk3247 n1088__vddio n1089__vddio 343.1e-3
rk3248 n1089__vddio n1090__vddio 52.73e-3
rk3249 n1090__vddio n1091__vddio 394.2e-3
rk3250 n1080__vddio n1081__vddio 3.1
rk3251 n1080__vddio n1084__vddio 3.1
rk3252 n1080__vddio n1087__vddio 3.1
rk3253 n1080__vddio n1090__vddio 3.1
rk3254 n619__vss n620__vss 55.24e-3
rk3255 n620__vss n621__vss 365.7e-3
rk3256 n621__vss n622__vss 298.6e-3
rk3257 n622__vss n623__vss 42.68e-3
rk3258 n623__vss n624__vss 365.7e-3
rk3259 n624__vss n625__vss 187.7e-3
rk3260 n625__vss n626__vss 264.6e-3
rk3261 n618__vss n619__vss 3.75
rk3262 n618__vss n622__vss 3.75
rk3263 n618__vss n625__vss 5.7692
rk3264 n706__i1__i14__net1 n769__i1__i14__net1 125e-3
rk3265 n708__i1__i14__net1 n770__i1__i14__net1 125e-3
rk3267 n22__shift n11__shift 45.0049
rk3268 n631__vss n632__vss 37.7533
rk3269 n151__vdd n153__vdd 70.25e-3
rk3270 n152__vdd n153__vdd 15.5
rk3271 n18__i5__i9__net21 n19__i5__i9__net21 15.9169
rk3272 n19__i5__i9__net21 n20__i5__i9__net21 37.8067
rk3273 n19__i5__i9__net21 n3__i5__i9__net21 22.7022
rk3275 n1891__chipdriverout n1893__chipdriverout 210.4e-3
rk3276 n1893__chipdriverout n1894__chipdriverout 155.3e-3
rk3277 n1894__chipdriverout n1895__chipdriverout 343.1e-3
rk3278 n1895__chipdriverout n1896__chipdriverout 226.6e-3
rk3279 n1896__chipdriverout n1897__chipdriverout 139.1e-3
rk3280 n1897__chipdriverout n1898__chipdriverout 362.5e-3
rk3281 n1898__chipdriverout n1899__chipdriverout 223.4e-3
rk3282 n1899__chipdriverout n1900__chipdriverout 142.4e-3
rk3283 n1900__chipdriverout n1901__chipdriverout 343.1e-3
rk3284 n1901__chipdriverout n1902__chipdriverout 239.6e-3
rk3285 n1902__chipdriverout n1903__chipdriverout 126.2e-3
rk3287 n1892__chipdriverout n1893__chipdriverout 3.1
rk3288 n1892__chipdriverout n1896__chipdriverout 3.1
rk3289 n1892__chipdriverout n1899__chipdriverout 3.1
rk3290 n1892__chipdriverout n1902__chipdriverout 3.1
rk3292 n1907__chipdriverout n1908__chipdriverout 12.55e-3
rk3293 n1908__chipdriverout n1909__chipdriverout 365.7e-3
rk3294 n1909__chipdriverout n1910__chipdriverout 226.6e-3
rk3295 n1910__chipdriverout n1911__chipdriverout 116.5e-3
rk3296 n1911__chipdriverout n1912__chipdriverout 365.7e-3
rk3297 n1912__chipdriverout n1913__chipdriverout 242.8e-3
rk3298 n1913__chipdriverout n1914__chipdriverout 119.7e-3
rk3300 n1906__chipdriverout n1907__chipdriverout 5.7692
rk3301 n1906__chipdriverout n1910__chipdriverout 3.75
rk3302 n1906__chipdriverout n1913__chipdriverout 3.75
rk3303 n714__i1__i14__net1 n773__i1__i14__net1 125e-3
rk3304 n716__i1__i14__net1 n774__i1__i14__net1 125e-3
rk3305 n156__vdd n157__vdd 320.2e-3
rk3306 n155__vdd n156__vdd 15.5
rk3307 n634__vss n635__vss 37.7549
rk3309 n1100__vddio n1102__vddio 30.13e-3
rk3310 n1102__vddio n1103__vddio 335.6e-3
rk3311 n1103__vddio n1104__vddio 343.1e-3
rk3312 n1104__vddio n1105__vddio 42.68e-3
rk3313 n1105__vddio n1106__vddio 321.2e-3
rk3314 n1106__vddio n1107__vddio 362.5e-3
rk3315 n1107__vddio n1108__vddio 40.17e-3
rk3316 n1108__vddio n1109__vddio 323.7e-3
rk3317 n1109__vddio n1110__vddio 343.1e-3
rk3318 n1110__vddio n1111__vddio 52.73e-3
rk3319 n1111__vddio n1112__vddio 394.2e-3
rk3320 n1101__vddio n1102__vddio 3.1
rk3321 n1101__vddio n1105__vddio 3.1
rk3322 n1101__vddio n1108__vddio 3.1
rk3323 n1101__vddio n1111__vddio 3.1
rk3324 n637__vss n638__vss 55.24e-3
rk3325 n638__vss n639__vss 365.7e-3
rk3326 n639__vss n640__vss 298.6e-3
rk3327 n640__vss n641__vss 42.68e-3
rk3328 n641__vss n642__vss 365.7e-3
rk3329 n642__vss n643__vss 187.7e-3
rk3330 n643__vss n644__vss 264.6e-3
rk3331 n636__vss n637__vss 3.75
rk3332 n636__vss n640__vss 3.75
rk3333 n636__vss n643__vss 5.7692
rk3334 n9__i5__i6__net32 n8__i5__i6__net32 31.2217
rk3335 n8__i5__i6__net32 n10__i5__i6__net32 75.2494
rk3336 n14__i5__i9__net21 n10__i5__i9__net21 119.4e-3
rk3337 n10__i5__i9__net21 n6__i5__i9__net21 119.4e-3
rk3338 n6__i5__i9__net21 i5__i9__net21 119.5e-3
rk3339 n16__i5__i9__net21 n12__i5__i9__net21 122.9e-3
rk3340 n12__i5__i9__net21 n8__i5__i9__net21 122.9e-3
rk3341 n8__i5__i9__net21 n5__i5__i9__net21 122.9e-3
rk3342 n700__vss n701__vss 4.9e-3
rk3343 n699__vss n700__vss 37.5
rk3344 n162__vdd n159__vdd 70.25e-3
rk3345 n161__vdd n162__vdd 15.5
rk3346 n10__i5__r1 n11__i5__r1 31.2117
rk3347 n11__i5__r1 n12__i5__r1 75.2117
rk3348 n4__i5__i6__i7__net4 n6__i5__i6__i7__net4 1.2154
rk3349 n6__i5__i6__i7__net4 n8__i5__i6__i7__net4 451.2e-3
rk3350 n8__i5__i6__i7__net4 n2__i5__i6__i7__net4 497.3e-3
rk3351 n5__i5__i6__i7__net4 n6__i5__i6__i7__net4 75
rk3352 n7__i5__i6__i7__net4 n8__i5__i6__i7__net4 31
rk3353 n20__shift n28__shift 1.3224
rk3354 n28__shift n18__shift 5.102e-3
rk3355 n8__i5__i6__net33 n9__i5__i6__net33 75.2457
rk3356 n9__i5__i6__net33 n11__i5__i6__net33 219e-3
rk3357 n11__i5__i6__net33 n13__i5__i6__net33 1.1197
rk3358 n13__i5__i6__net33 n14__i5__i6__net33 75.5378
rk3359 n10__i5__i6__net33 n11__i5__i6__net33 31
rk3360 n12__i5__i6__net33 n13__i5__i6__net33 31
rk3361 n21__i5__clk_buf n44__i5__clk_buf 22.5194
rk3362 n44__i5__clk_buf n45__i5__clk_buf 209.8e-3
rk3363 n45__i5__clk_buf n46__i5__clk_buf 122.6e-3
rk3364 n46__i5__clk_buf n47__i5__clk_buf 37.8139
rk3365 n45__i5__clk_buf n48__i5__clk_buf 37.8072
rk3366 n45__i5__clk_buf n49__i5__clk_buf 15.9139
rk3367 n46__i5__clk_buf n50__i5__clk_buf 15.9237
rk3368 n2__i5__i6__i4__net25 n3__i5__i6__i4__net25 323.3e-3
rk3369 i5__i6__i4__net25 n2__i5__i6__i4__net25 15.5
rk3370 i5__i6__i4__net21 n2__i5__i6__i4__net21 37.7516
rk3371 n3__i5__i6__net33 n15__i5__i6__net33 22.6237
rk3372 n8__i5__i8__net4 n9__i5__i8__net4 31.2664
rk3373 n9__i5__i8__net4 n10__i5__i8__net4 289.5e-3
rk3374 n10__i5__i8__net4 n11__i5__i8__net4 75.2485
rk3375 n9__i5__i8__net4 n12__i5__i8__net4 34.67e-3
rk3376 n12__i5__i8__net4 n13__i5__i8__net4 75.0632
rk3377 n10__i5__i8__net4 n14__i5__i8__net4 31.3077
rk3378 n5__i5__i6__i4__net25 n6__i5__i6__i4__net25 350.8e-3
rk3379 n4__i5__i6__i4__net25 n5__i5__i6__i4__net25 15.5
rk3380 n3__i5__i6__i4__net21 n5__i5__i6__i4__net21 4.9e-3
rk3381 n4__i5__i6__i4__net21 n5__i5__i6__i4__net21 37.5
rk3382 n20__i5__i6__net31 n29__i5__i6__net31 500e-3
rk3383 n31__i5__clk_buf n51__i5__clk_buf 500e-3
rk3384 n2__i5__i8__i9__net25 n3__i5__i8__i9__net25 323.3e-3
rk3385 i5__i8__i9__net25 n2__i5__i8__i9__net25 15.5
rk3386 i5__i8__i9__net21 n2__i5__i8__i9__net21 37.7516
rk3387 n8__i5__i6__i4__net25 n9__i5__i6__i4__net25 350.8e-3
rk3388 n7__i5__i6__i4__net25 n8__i5__i6__i4__net25 15.5
rk3389 n6__i5__i6__i4__net21 n8__i5__i6__i4__net21 4.9e-3
rk3390 n7__i5__i6__i4__net21 n8__i5__i6__i4__net21 37.5
rk3391 n9__i5__i8__net1 n3__i5__i8__net1 22.558
rk3393 n1174__vddio n1176__vddio 30.13e-3
rk3394 n1176__vddio n1177__vddio 335.6e-3
rk3395 n1177__vddio n1178__vddio 343.1e-3
rk3396 n1178__vddio n1179__vddio 42.68e-3
rk3397 n1179__vddio n1180__vddio 321.2e-3
rk3398 n1180__vddio n1181__vddio 362.5e-3
rk3399 n1181__vddio n1182__vddio 40.17e-3
rk3400 n1182__vddio n1183__vddio 323.7e-3
rk3401 n1183__vddio n1184__vddio 343.1e-3
rk3402 n1184__vddio n1185__vddio 52.73e-3
rk3403 n1185__vddio n1186__vddio 394.2e-3
rk3404 n1175__vddio n1176__vddio 3.1
rk3405 n1175__vddio n1179__vddio 3.1
rk3406 n1175__vddio n1182__vddio 3.1
rk3407 n1175__vddio n1185__vddio 3.1
rk3408 n704__vss n705__vss 55.24e-3
rk3409 n705__vss n706__vss 365.7e-3
rk3410 n706__vss n707__vss 298.6e-3
rk3411 n707__vss n708__vss 42.68e-3
rk3412 n708__vss n709__vss 365.7e-3
rk3413 n709__vss n710__vss 187.7e-3
rk3414 n710__vss n711__vss 264.6e-3
rk3415 n703__vss n704__vss 3.75
rk3416 n703__vss n707__vss 3.75
rk3417 n703__vss n710__vss 5.7692
rk3418 n5__i5__i8__i9__net25 n6__i5__i8__i9__net25 350.8e-3
rk3419 n4__i5__i8__i9__net25 n5__i5__i8__i9__net25 15.5
rk3420 n3__i5__i8__i9__net21 n5__i5__i8__i9__net21 4.9e-3
rk3421 n4__i5__i8__i9__net21 n5__i5__i8__i9__net21 37.5
rk3422 n3__i5__i8__net4 n15__i5__i8__net4 500e-3
rk3423 n2__i5__i6__i4__net24 n3__i5__i6__i4__net24 323.3e-3
rk3424 i5__i6__i4__net24 n2__i5__i6__i4__net24 15.5
rk3425 i5__i6__i4__net23 n2__i5__i6__i4__net23 37.7516
rk3426 i1__net2 n61__i1__net2 125e-3
rk3427 n3__i1__net2 n62__i1__net2 125e-3
rk3428 n34__i5__clk_buf n56__i5__clk_buf 500e-3
rk3430 n793__i1__i14__net1 n794__i1__i14__net1 12.55e-3
rk3431 n794__i1__i14__net1 n795__i1__i14__net1 365.7e-3
rk3432 n795__i1__i14__net1 n796__i1__i14__net1 226.6e-3
rk3433 n796__i1__i14__net1 n797__i1__i14__net1 116.5e-3
rk3434 n797__i1__i14__net1 n798__i1__i14__net1 365.7e-3
rk3435 n798__i1__i14__net1 n799__i1__i14__net1 242.8e-3
rk3436 n799__i1__i14__net1 n800__i1__i14__net1 119.7e-3
rk3438 n792__i1__i14__net1 n793__i1__i14__net1 5.7692
rk3439 n792__i1__i14__net1 n796__i1__i14__net1 3.75
rk3440 n792__i1__i14__net1 n799__i1__i14__net1 3.75
rk3442 n803__i1__i14__net1 n805__i1__i14__net1 210.4e-3
rk3443 n805__i1__i14__net1 n806__i1__i14__net1 155.3e-3
rk3444 n806__i1__i14__net1 n807__i1__i14__net1 343.1e-3
rk3445 n807__i1__i14__net1 n808__i1__i14__net1 226.6e-3
rk3446 n808__i1__i14__net1 n809__i1__i14__net1 139.1e-3
rk3447 n809__i1__i14__net1 n810__i1__i14__net1 362.5e-3
rk3448 n810__i1__i14__net1 n811__i1__i14__net1 223.4e-3
rk3449 n811__i1__i14__net1 n812__i1__i14__net1 142.4e-3
rk3450 n812__i1__i14__net1 n813__i1__i14__net1 343.1e-3
rk3451 n813__i1__i14__net1 n814__i1__i14__net1 239.6e-3
rk3452 n814__i1__i14__net1 n815__i1__i14__net1 126.2e-3
rk3454 n804__i1__i14__net1 n805__i1__i14__net1 3.1
rk3455 n804__i1__i14__net1 n808__i1__i14__net1 3.1
rk3456 n804__i1__i14__net1 n811__i1__i14__net1 3.1
rk3457 n804__i1__i14__net1 n814__i1__i14__net1 3.1
rk3458 n8__i5__i6__i4__net22 n9__i5__i6__i4__net22 15.9814
rk3459 n9__i5__i6__i4__net22 n10__i5__i6__i4__net22 37.8249
rk3460 n9__i5__i6__i4__net22 n3__i5__i6__i4__net22 22.9156
rk3461 n8__i5__i8__i9__net25 n9__i5__i8__i9__net25 350.8e-3
rk3462 n7__i5__i8__i9__net25 n8__i5__i8__i9__net25 15.5
rk3463 n6__i5__i8__i9__net21 n8__i5__i8__i9__net21 4.9e-3
rk3464 n7__i5__i8__i9__net21 n8__i5__i8__i9__net21 37.5
rk3465 n6__i1__net2 n69__i1__net2 125e-3
rk3466 n8__i1__net2 n70__i1__net2 125e-3
rk3467 n5__i5__i6__i4__net24 n6__i5__i6__i4__net24 350.8e-3
rk3468 n4__i5__i6__i4__net24 n5__i5__i6__i4__net24 15.5
rk3469 n3__i5__i6__i4__net23 n5__i5__i6__i4__net23 4.9e-3
rk3470 n4__i5__i6__i4__net23 n5__i5__i6__i4__net23 37.5
rk3472 n1201__vddio n1203__vddio 30.13e-3
rk3473 n1203__vddio n1204__vddio 335.6e-3
rk3474 n1204__vddio n1205__vddio 343.1e-3
rk3475 n1205__vddio n1206__vddio 42.68e-3
rk3476 n1206__vddio n1207__vddio 321.2e-3
rk3477 n1207__vddio n1208__vddio 362.5e-3
rk3478 n1208__vddio n1209__vddio 40.17e-3
rk3479 n1209__vddio n1210__vddio 323.7e-3
rk3480 n1210__vddio n1211__vddio 343.1e-3
rk3481 n1211__vddio n1212__vddio 52.73e-3
rk3482 n1212__vddio n1213__vddio 394.2e-3
rk3483 n1202__vddio n1203__vddio 3.1
rk3484 n1202__vddio n1206__vddio 3.1
rk3485 n1202__vddio n1209__vddio 3.1
rk3486 n1202__vddio n1212__vddio 3.1
rk3487 n717__vss n718__vss 55.24e-3
rk3488 n718__vss n719__vss 365.7e-3
rk3489 n719__vss n720__vss 298.6e-3
rk3490 n720__vss n721__vss 42.68e-3
rk3491 n721__vss n722__vss 365.7e-3
rk3492 n722__vss n723__vss 187.7e-3
rk3493 n723__vss n724__vss 264.6e-3
rk3494 n716__vss n717__vss 3.75
rk3495 n716__vss n720__vss 3.75
rk3496 n716__vss n723__vss 5.7692
rk3498 n39__i5__clk_buf n58__i5__clk_buf 500e-3
rk3499 n2__i5__i8__i9__net24 n3__i5__i8__i9__net24 323.3e-3
rk3500 i5__i8__i9__net24 n2__i5__i8__i9__net24 15.5
rk3501 i5__i8__i9__net23 n2__i5__i8__i9__net23 37.7516
rk3502 n9__i1__net2 n77__i1__net2 125e-3
rk3503 n11__i1__net2 n78__i1__net2 125e-3
rk3504 n8__i5__i6__i4__net24 n9__i5__i6__i4__net24 350.8e-3
rk3505 n7__i5__i6__i4__net24 n8__i5__i6__i4__net24 15.5
rk3506 n6__i5__i6__i4__net23 n8__i5__i6__i4__net23 4.9e-3
rk3507 n7__i5__i6__i4__net23 n8__i5__i6__i4__net23 37.5
rk3509 n832__i1__i14__net1 n833__i1__i14__net1 12.55e-3
rk3510 n833__i1__i14__net1 n834__i1__i14__net1 365.7e-3
rk3511 n834__i1__i14__net1 n835__i1__i14__net1 226.6e-3
rk3512 n835__i1__i14__net1 n836__i1__i14__net1 116.5e-3
rk3513 n836__i1__i14__net1 n837__i1__i14__net1 365.7e-3
rk3514 n837__i1__i14__net1 n838__i1__i14__net1 242.8e-3
rk3515 n838__i1__i14__net1 n839__i1__i14__net1 119.7e-3
rk3517 n831__i1__i14__net1 n832__i1__i14__net1 5.7692
rk3518 n831__i1__i14__net1 n835__i1__i14__net1 3.75
rk3519 n831__i1__i14__net1 n838__i1__i14__net1 3.75
rk3521 n842__i1__i14__net1 n844__i1__i14__net1 210.4e-3
rk3522 n844__i1__i14__net1 n845__i1__i14__net1 155.3e-3
rk3523 n845__i1__i14__net1 n846__i1__i14__net1 343.1e-3
rk3524 n846__i1__i14__net1 n847__i1__i14__net1 226.6e-3
rk3525 n847__i1__i14__net1 n848__i1__i14__net1 139.1e-3
rk3526 n848__i1__i14__net1 n849__i1__i14__net1 362.5e-3
rk3527 n849__i1__i14__net1 n850__i1__i14__net1 223.4e-3
rk3528 n850__i1__i14__net1 n851__i1__i14__net1 142.4e-3
rk3529 n851__i1__i14__net1 n852__i1__i14__net1 343.1e-3
rk3530 n852__i1__i14__net1 n853__i1__i14__net1 239.6e-3
rk3531 n853__i1__i14__net1 n854__i1__i14__net1 126.2e-3
rk3533 n843__i1__i14__net1 n844__i1__i14__net1 3.1
rk3534 n843__i1__i14__net1 n847__i1__i14__net1 3.1
rk3535 n843__i1__i14__net1 n850__i1__i14__net1 3.1
rk3536 n843__i1__i14__net1 n853__i1__i14__net1 3.1
rk3537 n8__i5__i8__i9__net22 n9__i5__i8__i9__net22 15.9814
rk3538 n9__i5__i8__i9__net22 n10__i5__i8__i9__net22 37.8249
rk3539 n9__i5__i8__i9__net22 n3__i5__i8__i9__net22 22.9156
rk3543 n5__i5__i8__i9__net24 n6__i5__i8__i9__net24 350.8e-3
rk3544 n4__i5__i8__i9__net24 n5__i5__i8__i9__net24 15.5
rk3545 n3__i5__i8__i9__net23 n5__i5__i8__i9__net23 4.9e-3
rk3546 n4__i5__i8__i9__net23 n5__i5__i8__i9__net23 37.5
rk3547 n730__vss n731__vss 55.24e-3
rk3548 n731__vss n732__vss 365.7e-3
rk3549 n732__vss n733__vss 298.6e-3
rk3550 n733__vss n734__vss 42.68e-3
rk3551 n734__vss n735__vss 365.7e-3
rk3552 n735__vss n736__vss 187.7e-3
rk3553 n736__vss n737__vss 264.6e-3
rk3554 n729__vss n730__vss 3.75
rk3555 n729__vss n733__vss 3.75
rk3556 n729__vss n736__vss 5.7692
rk3558 n1222__vddio n1224__vddio 30.13e-3
rk3559 n1224__vddio n1225__vddio 335.6e-3
rk3560 n1225__vddio n1226__vddio 343.1e-3
rk3561 n1226__vddio n1227__vddio 42.68e-3
rk3562 n1227__vddio n1228__vddio 321.2e-3
rk3563 n1228__vddio n1229__vddio 362.5e-3
rk3564 n1229__vddio n1230__vddio 40.17e-3
rk3565 n1230__vddio n1231__vddio 323.7e-3
rk3566 n1231__vddio n1232__vddio 343.1e-3
rk3567 n1232__vddio n1233__vddio 52.73e-3
rk3568 n1233__vddio n1234__vddio 394.2e-3
rk3569 n1223__vddio n1224__vddio 3.1
rk3570 n1223__vddio n1227__vddio 3.1
rk3571 n1223__vddio n1230__vddio 3.1
rk3572 n1223__vddio n1233__vddio 3.1
rk3574 n42__i5__clk_buf n63__i5__clk_buf 500e-3
rk3575 n18__i1__net2 n89__i1__net2 125e-3
rk3576 n20__i1__net2 n90__i1__net2 125e-3
rk3577 n9__i5__i8__i9__net24 n7__i5__i8__i9__net24 100.8e-3
rk3578 n8__i5__i8__i9__net24 n9__i5__i8__i9__net24 15.5
rk3579 n6__i5__i8__i9__net23 n9__i5__i8__i9__net23 4.9e-3
rk3580 n8__i5__i8__i9__net23 n9__i5__i8__i9__net23 37.5
rk3582 n871__i1__i14__net1 n872__i1__i14__net1 12.55e-3
rk3583 n872__i1__i14__net1 n873__i1__i14__net1 365.7e-3
rk3584 n873__i1__i14__net1 n874__i1__i14__net1 226.6e-3
rk3585 n874__i1__i14__net1 n875__i1__i14__net1 116.5e-3
rk3586 n875__i1__i14__net1 n876__i1__i14__net1 365.7e-3
rk3587 n876__i1__i14__net1 n877__i1__i14__net1 242.8e-3
rk3588 n877__i1__i14__net1 n878__i1__i14__net1 119.7e-3
rk3590 n870__i1__i14__net1 n871__i1__i14__net1 5.7692
rk3591 n870__i1__i14__net1 n874__i1__i14__net1 3.75
rk3592 n870__i1__i14__net1 n877__i1__i14__net1 3.75
rk3594 n881__i1__i14__net1 n883__i1__i14__net1 212.2e-3
rk3595 n883__i1__i14__net1 n884__i1__i14__net1 157.2e-3
rk3596 n884__i1__i14__net1 n885__i1__i14__net1 346.7e-3
rk3597 n885__i1__i14__net1 n886__i1__i14__net1 228.4e-3
rk3598 n886__i1__i14__net1 n887__i1__i14__net1 141e-3
rk3599 n887__i1__i14__net1 n888__i1__i14__net1 366.1e-3
rk3600 n888__i1__i14__net1 n889__i1__i14__net1 225.2e-3
rk3601 n889__i1__i14__net1 n890__i1__i14__net1 144.2e-3
rk3602 n890__i1__i14__net1 n891__i1__i14__net1 346.7e-3
rk3603 n891__i1__i14__net1 n892__i1__i14__net1 241.4e-3
rk3604 n892__i1__i14__net1 n893__i1__i14__net1 128e-3
rk3606 n882__i1__i14__net1 n883__i1__i14__net1 3.1
rk3607 n882__i1__i14__net1 n886__i1__i14__net1 3.1
rk3608 n882__i1__i14__net1 n889__i1__i14__net1 3.1
rk3609 n882__i1__i14__net1 n892__i1__i14__net1 3.1
rk3610 i5__i6__net34 n2__i5__i6__net34 19.0545
rk3611 n2__i5__i6__net34 n3__i5__i6__net34 300.1e-3
rk3612 n3__i5__i6__net34 n4__i5__i6__net34 420.4e-3
rk3613 n4__i5__i6__net34 n5__i5__i6__net34 37.828
rk3614 n3__i5__i6__net34 n6__i5__i6__net34 19.0309
rk3615 n4__i5__i6__net34 n7__i5__i6__net34 15.8422
rk3616 n22__i1__net2 n97__i1__net2 125e-3
rk3617 n24__i1__net2 n98__i1__net2 125e-3
rk3618 n49__reset n54__reset 250e-3
rk3619 n751__vss n748__vss 55.24e-3
rk3620 n748__vss n747__vss 365.7e-3
rk3621 n747__vss n752__vss 298.6e-3
rk3622 n752__vss n744__vss 42.68e-3
rk3623 n744__vss n743__vss 365.7e-3
rk3624 n743__vss n753__vss 187.7e-3
rk3625 n753__vss n754__vss 264.6e-3
rk3626 n750__vss n751__vss 3.75
rk3627 n750__vss n752__vss 3.75
rk3628 n750__vss n753__vss 5.7692
rk3630 n1243__vddio n1258__vddio 30.13e-3
rk3631 n1258__vddio n1244__vddio 335.6e-3
rk3632 n1244__vddio n1247__vddio 343.1e-3
rk3633 n1247__vddio n1259__vddio 42.68e-3
rk3634 n1259__vddio n1248__vddio 321.2e-3
rk3635 n1248__vddio n1251__vddio 362.5e-3
rk3636 n1251__vddio n1260__vddio 40.17e-3
rk3637 n1260__vddio n1252__vddio 323.7e-3
rk3638 n1252__vddio n1255__vddio 343.1e-3
rk3639 n1255__vddio n1261__vddio 52.73e-3
rk3640 n1261__vddio n1262__vddio 394.2e-3
rk3641 n1257__vddio n1258__vddio 3.1
rk3642 n1257__vddio n1259__vddio 3.1
rk3643 n1257__vddio n1260__vddio 3.1
rk3644 n1257__vddio n1261__vddio 3.1
rk3646 n35__shift n24__shift 45.0049
rk3647 n26__i1__net2 n109__i1__net2 125e-3
rk3648 n28__i1__net2 n110__i1__net2 125e-3
rk3650 n910__i1__i14__net1 n911__i1__i14__net1 12.55e-3
rk3651 n911__i1__i14__net1 n912__i1__i14__net1 365.7e-3
rk3652 n912__i1__i14__net1 n913__i1__i14__net1 226.6e-3
rk3653 n913__i1__i14__net1 n914__i1__i14__net1 116.5e-3
rk3654 n914__i1__i14__net1 n915__i1__i14__net1 365.7e-3
rk3655 n915__i1__i14__net1 n916__i1__i14__net1 242.8e-3
rk3656 n916__i1__i14__net1 n917__i1__i14__net1 119.7e-3
rk3658 n909__i1__i14__net1 n910__i1__i14__net1 5.7692
rk3659 n909__i1__i14__net1 n913__i1__i14__net1 3.75
rk3660 n909__i1__i14__net1 n916__i1__i14__net1 3.75
rk3662 n920__i1__i14__net1 n922__i1__i14__net1 212.2e-3
rk3663 n922__i1__i14__net1 n923__i1__i14__net1 157.2e-3
rk3664 n923__i1__i14__net1 n924__i1__i14__net1 346.7e-3
rk3665 n924__i1__i14__net1 n925__i1__i14__net1 228.4e-3
rk3666 n925__i1__i14__net1 n926__i1__i14__net1 141e-3
rk3667 n926__i1__i14__net1 n927__i1__i14__net1 366.1e-3
rk3668 n927__i1__i14__net1 n928__i1__i14__net1 225.2e-3
rk3669 n928__i1__i14__net1 n929__i1__i14__net1 144.2e-3
rk3670 n929__i1__i14__net1 n930__i1__i14__net1 346.7e-3
rk3671 n930__i1__i14__net1 n931__i1__i14__net1 241.4e-3
rk3672 n931__i1__i14__net1 n932__i1__i14__net1 128e-3
rk3674 n921__i1__i14__net1 n922__i1__i14__net1 3.1
rk3675 n921__i1__i14__net1 n925__i1__i14__net1 3.1
rk3676 n921__i1__i14__net1 n928__i1__i14__net1 3.1
rk3677 n921__i1__i14__net1 n931__i1__i14__net1 3.1
rk3680 n9__i5__i6__net34 n8__i5__i6__net34 31.2217
rk3681 n8__i5__i6__net34 n10__i5__i6__net34 75.2494
rk3683 n1264__vddio n1266__vddio 30.13e-3
rk3684 n1266__vddio n1267__vddio 335.6e-3
rk3685 n1267__vddio n1268__vddio 343.1e-3
rk3686 n1268__vddio n1269__vddio 42.68e-3
rk3687 n1269__vddio n1270__vddio 321.2e-3
rk3688 n1270__vddio n1271__vddio 362.5e-3
rk3689 n1271__vddio n1272__vddio 40.17e-3
rk3690 n1272__vddio n1273__vddio 323.7e-3
rk3691 n1273__vddio n1274__vddio 343.1e-3
rk3692 n1274__vddio n1275__vddio 52.73e-3
rk3693 n1275__vddio n1276__vddio 394.2e-3
rk3694 n1265__vddio n1266__vddio 3.1
rk3695 n1265__vddio n1269__vddio 3.1
rk3696 n1265__vddio n1272__vddio 3.1
rk3697 n1265__vddio n1275__vddio 3.1
rk3698 n756__vss n757__vss 55.24e-3
rk3699 n757__vss n758__vss 365.7e-3
rk3700 n758__vss n759__vss 298.6e-3
rk3701 n759__vss n760__vss 42.68e-3
rk3702 n760__vss n761__vss 365.7e-3
rk3703 n761__vss n762__vss 187.7e-3
rk3704 n762__vss n763__vss 264.6e-3
rk3705 n755__vss n756__vss 3.75
rk3706 n755__vss n759__vss 3.75
rk3707 n755__vss n762__vss 5.7692
rk3710 n17__i5__i8__net2 n20__i5__i8__net2 428.8e-3
rk3711 n20__i5__i8__net2 n21__i5__i8__net2 131.7e-3
rk3712 n21__i5__i8__net2 n22__i5__i8__net2 87.73e-3
rk3713 n22__i5__i8__net2 n23__i5__i8__net2 204e-3
rk3714 n23__i5__i8__net2 n24__i5__i8__net2 420.4e-3
rk3715 n24__i5__i8__net2 n25__i5__i8__net2 37.828
rk3716 n20__i5__i8__net2 n4__i5__i8__net2 22.7212
rk3717 n21__i5__i8__net2 n26__i5__i8__net2 19.0331
rk3718 n22__i5__i8__net2 n27__i5__i8__net2 637.7e-3
rk3719 n23__i5__i8__net2 n28__i5__i8__net2 19.0331
rk3720 n24__i5__i8__net2 n29__i5__i8__net2 15.8422
rk3722 n949__i1__i14__net1 n950__i1__i14__net1 12.55e-3
rk3723 n950__i1__i14__net1 n951__i1__i14__net1 365.7e-3
rk3724 n951__i1__i14__net1 n952__i1__i14__net1 226.6e-3
rk3725 n952__i1__i14__net1 n953__i1__i14__net1 116.5e-3
rk3726 n953__i1__i14__net1 n954__i1__i14__net1 365.7e-3
rk3727 n954__i1__i14__net1 n955__i1__i14__net1 242.8e-3
rk3728 n955__i1__i14__net1 n956__i1__i14__net1 119.7e-3
rk3730 n948__i1__i14__net1 n949__i1__i14__net1 5.7692
rk3731 n948__i1__i14__net1 n952__i1__i14__net1 3.75
rk3732 n948__i1__i14__net1 n955__i1__i14__net1 3.75
rk3734 n959__i1__i14__net1 n961__i1__i14__net1 210.4e-3
rk3735 n961__i1__i14__net1 n962__i1__i14__net1 155.3e-3
rk3736 n962__i1__i14__net1 n963__i1__i14__net1 343.1e-3
rk3737 n963__i1__i14__net1 n964__i1__i14__net1 226.6e-3
rk3738 n964__i1__i14__net1 n965__i1__i14__net1 139.1e-3
rk3739 n965__i1__i14__net1 n966__i1__i14__net1 362.5e-3
rk3740 n966__i1__i14__net1 n967__i1__i14__net1 223.4e-3
rk3741 n967__i1__i14__net1 n968__i1__i14__net1 142.4e-3
rk3742 n968__i1__i14__net1 n969__i1__i14__net1 343.1e-3
rk3743 n969__i1__i14__net1 n970__i1__i14__net1 239.6e-3
rk3744 n970__i1__i14__net1 n971__i1__i14__net1 126.2e-3
rk3746 n960__i1__i14__net1 n961__i1__i14__net1 3.1
rk3747 n960__i1__i14__net1 n964__i1__i14__net1 3.1
rk3748 n960__i1__i14__net1 n967__i1__i14__net1 3.1
rk3749 n960__i1__i14__net1 n970__i1__i14__net1 3.1
rk3750 n38__i1__net2 n129__i1__net2 125e-3
rk3751 n40__i1__net2 n130__i1__net2 125e-3
rk3752 n11__i5__r0 n12__i5__r0 31.2117
rk3753 n12__i5__r0 n13__i5__r0 75.2117
rk3754 n4__i5__i6__i8__net4 n6__i5__i6__i8__net4 1.2154
rk3755 n6__i5__i6__i8__net4 n8__i5__i6__i8__net4 451.2e-3
rk3756 n8__i5__i6__i8__net4 n2__i5__i6__i8__net4 497.3e-3
rk3757 n5__i5__i6__i8__net4 n6__i5__i6__i8__net4 75
rk3758 n7__i5__i6__i8__net4 n8__i5__i6__i8__net4 31
rk3759 n33__shift n38__shift 1.3224
rk3760 n38__shift n31__shift 5.102e-3
rk3762 n1295__vddio n1297__vddio 30.13e-3
rk3763 n1297__vddio n1298__vddio 335.6e-3
rk3764 n1298__vddio n1299__vddio 343.1e-3
rk3765 n1299__vddio n1300__vddio 42.68e-3
rk3766 n1300__vddio n1301__vddio 321.2e-3
rk3767 n1301__vddio n1302__vddio 362.5e-3
rk3768 n1302__vddio n1303__vddio 40.17e-3
rk3769 n1303__vddio n1304__vddio 323.7e-3
rk3770 n1304__vddio n1305__vddio 343.1e-3
rk3771 n1305__vddio n1306__vddio 52.73e-3
rk3772 n1306__vddio n1307__vddio 394.2e-3
rk3773 n1296__vddio n1297__vddio 3.1
rk3774 n1296__vddio n1300__vddio 3.1
rk3775 n1296__vddio n1303__vddio 3.1
rk3776 n1296__vddio n1306__vddio 3.1
rk3777 n769__vss n770__vss 55.24e-3
rk3778 n770__vss n771__vss 365.7e-3
rk3779 n771__vss n772__vss 298.6e-3
rk3780 n772__vss n773__vss 42.68e-3
rk3781 n773__vss n774__vss 365.7e-3
rk3782 n774__vss n775__vss 187.7e-3
rk3783 n775__vss n776__vss 264.6e-3
rk3784 n768__vss n769__vss 3.75
rk3785 n768__vss n772__vss 3.75
rk3786 n768__vss n775__vss 5.7692
rk3787 n8__i5__i6__net35 n9__i5__i6__net35 75.2457
rk3788 n9__i5__i6__net35 n11__i5__i6__net35 219e-3
rk3789 n11__i5__i6__net35 n13__i5__i6__net35 1.1197
rk3790 n13__i5__i6__net35 n14__i5__i6__net35 75.5378
rk3791 n10__i5__i6__net35 n11__i5__i6__net35 31
rk3792 n12__i5__i6__net35 n13__i5__i6__net35 31
rk3793 n42__i1__net2 n141__i1__net2 125e-3
rk3794 n44__i1__net2 n142__i1__net2 125e-3
rk3795 n18__i5__i8__net1 n19__i5__i8__net1 31.2678
rk3796 n19__i5__i8__net1 n20__i5__i8__net1 291.7e-3
rk3797 n20__i5__i8__net1 n21__i5__i8__net1 75.2422
rk3798 n19__i5__i8__net1 n22__i5__i8__net1 75.1768
rk3799 n20__i5__i8__net1 n23__i5__i8__net1 31.3039
rk3801 n988__i1__i14__net1 n989__i1__i14__net1 12.55e-3
rk3802 n989__i1__i14__net1 n990__i1__i14__net1 365.7e-3
rk3803 n990__i1__i14__net1 n991__i1__i14__net1 226.6e-3
rk3804 n991__i1__i14__net1 n992__i1__i14__net1 116.5e-3
rk3805 n992__i1__i14__net1 n993__i1__i14__net1 365.7e-3
rk3806 n993__i1__i14__net1 n994__i1__i14__net1 242.8e-3
rk3807 n994__i1__i14__net1 n995__i1__i14__net1 119.7e-3
rk3809 n987__i1__i14__net1 n988__i1__i14__net1 5.7692
rk3810 n987__i1__i14__net1 n991__i1__i14__net1 3.75
rk3811 n987__i1__i14__net1 n994__i1__i14__net1 3.75
rk3813 n998__i1__i14__net1 n1000__i1__i14__net1 210.4e-3
rk3814 n1000__i1__i14__net1 n1001__i1__i14__net1 155.3e-3
rk3815 n1001__i1__i14__net1 n1002__i1__i14__net1 343.1e-3
rk3816 n1002__i1__i14__net1 n1003__i1__i14__net1 226.6e-3
rk3817 n1003__i1__i14__net1 n1004__i1__i14__net1 139.1e-3
rk3818 n1004__i1__i14__net1 n1005__i1__i14__net1 362.5e-3
rk3819 n1005__i1__i14__net1 n1006__i1__i14__net1 223.4e-3
rk3820 n1006__i1__i14__net1 n1007__i1__i14__net1 142.4e-3
rk3821 n1007__i1__i14__net1 n1008__i1__i14__net1 343.1e-3
rk3822 n1008__i1__i14__net1 n1009__i1__i14__net1 239.6e-3
rk3823 n1009__i1__i14__net1 n1010__i1__i14__net1 126.2e-3
rk3825 n999__i1__i14__net1 n1000__i1__i14__net1 3.1
rk3826 n999__i1__i14__net1 n1003__i1__i14__net1 3.1
rk3827 n999__i1__i14__net1 n1006__i1__i14__net1 3.1
rk3828 n999__i1__i14__net1 n1009__i1__i14__net1 3.1
rk3829 n2__i5__i6__i5__net25 n3__i5__i6__i5__net25 323.3e-3
rk3830 i5__i6__i5__net25 n2__i5__i6__i5__net25 15.5
rk3831 i5__i6__i5__net21 n2__i5__i6__i5__net21 37.7516
rk3832 n2__i5__i8__i10__net25 n3__i5__i8__i10__net25 323.3e-3
rk3833 i5__i8__i10__net25 n2__i5__i8__i10__net25 15.5
rk3834 i5__i8__i10__net21 n2__i5__i8__i10__net21 37.7516
rk3835 n46__i1__net2 n149__i1__net2 125e-3
rk3836 n48__i1__net2 n150__i1__net2 125e-3
rk3837 n3__i5__i6__net35 n15__i5__i6__net35 22.6237
rk3838 n782__vss n783__vss 55.24e-3
rk3839 n783__vss n784__vss 365.7e-3
rk3840 n784__vss n785__vss 298.6e-3
rk3841 n785__vss n786__vss 42.68e-3
rk3842 n786__vss n787__vss 365.7e-3
rk3843 n787__vss n788__vss 187.7e-3
rk3844 n788__vss n789__vss 264.6e-3
rk3845 n781__vss n782__vss 3.75
rk3846 n781__vss n785__vss 3.75
rk3847 n781__vss n788__vss 5.7692
rk3849 n1316__vddio n1318__vddio 30.13e-3
rk3850 n1318__vddio n1319__vddio 335.6e-3
rk3851 n1319__vddio n1320__vddio 343.1e-3
rk3852 n1320__vddio n1321__vddio 42.68e-3
rk3853 n1321__vddio n1322__vddio 321.2e-3
rk3854 n1322__vddio n1323__vddio 362.5e-3
rk3855 n1323__vddio n1324__vddio 40.17e-3
rk3856 n1324__vddio n1325__vddio 323.7e-3
rk3857 n1325__vddio n1326__vddio 343.1e-3
rk3858 n1326__vddio n1327__vddio 52.73e-3
rk3859 n1327__vddio n1328__vddio 394.2e-3
rk3860 n1317__vddio n1318__vddio 3.1
rk3861 n1317__vddio n1321__vddio 3.1
rk3862 n1317__vddio n1324__vddio 3.1
rk3863 n1317__vddio n1327__vddio 3.1
rk3864 n3__i5__i8__net5 n8__i5__i8__net5 22.7766
rk3865 n5__i5__i6__i5__net25 n6__i5__i6__i5__net25 350.8e-3
rk3866 n4__i5__i6__i5__net25 n5__i5__i6__i5__net25 15.5
rk3867 n3__i5__i6__i5__net21 n5__i5__i6__i5__net21 4.9e-3
rk3868 n4__i5__i6__i5__net21 n5__i5__i6__i5__net21 37.5
rk3869 n50__i1__net2 n157__i1__net2 125e-3
rk3870 n52__i1__net2 n158__i1__net2 125e-3
rk3871 n5__i5__i8__i10__net25 n6__i5__i8__i10__net25 350.8e-3
rk3872 n4__i5__i8__i10__net25 n5__i5__i8__i10__net25 15.5
rk3873 n3__i5__i8__i10__net21 n5__i5__i8__i10__net21 4.9e-3
rk3874 n4__i5__i8__i10__net21 n5__i5__i8__i10__net21 37.5
rk3875 n34__i5__i6__net31 n41__i5__i6__net31 500e-3
rk3876 n13__i5__i8__net1 n26__i5__i8__net1 500e-3
rk3877 n55__i5__clk_buf n65__i5__clk_buf 500e-3
rk3879 n1026__i1__i14__net1 n1028__i1__i14__net1 210.4e-3
rk3880 n1028__i1__i14__net1 n1029__i1__i14__net1 155.3e-3
rk3881 n1029__i1__i14__net1 n1030__i1__i14__net1 343.1e-3
rk3882 n1030__i1__i14__net1 n1031__i1__i14__net1 226.6e-3
rk3883 n1031__i1__i14__net1 n1032__i1__i14__net1 139.1e-3
rk3884 n1032__i1__i14__net1 n1033__i1__i14__net1 362.5e-3
rk3885 n1033__i1__i14__net1 n1034__i1__i14__net1 223.4e-3
rk3886 n1034__i1__i14__net1 n1035__i1__i14__net1 142.4e-3
rk3887 n1035__i1__i14__net1 n1036__i1__i14__net1 343.1e-3
rk3888 n1036__i1__i14__net1 n1037__i1__i14__net1 239.6e-3
rk3889 n1037__i1__i14__net1 n1038__i1__i14__net1 126.2e-3
rk3891 n1027__i1__i14__net1 n1028__i1__i14__net1 3.1
rk3892 n1027__i1__i14__net1 n1031__i1__i14__net1 3.1
rk3893 n1027__i1__i14__net1 n1034__i1__i14__net1 3.1
rk3894 n1027__i1__i14__net1 n1037__i1__i14__net1 3.1
rk3896 n1042__i1__i14__net1 n1043__i1__i14__net1 12.55e-3
rk3897 n1043__i1__i14__net1 n1044__i1__i14__net1 365.7e-3
rk3898 n1044__i1__i14__net1 n1045__i1__i14__net1 226.6e-3
rk3899 n1045__i1__i14__net1 n1046__i1__i14__net1 116.5e-3
rk3900 n1046__i1__i14__net1 n1047__i1__i14__net1 365.7e-3
rk3901 n1047__i1__i14__net1 n1048__i1__i14__net1 242.8e-3
rk3902 n1048__i1__i14__net1 n1049__i1__i14__net1 119.7e-3
rk3904 n1041__i1__i14__net1 n1042__i1__i14__net1 5.7692
rk3905 n1041__i1__i14__net1 n1045__i1__i14__net1 3.75
rk3906 n1041__i1__i14__net1 n1048__i1__i14__net1 3.75
rk3907 n12__i5__i8__net2 n33__i5__i8__net2 500e-3
rk3910 n9__i5__i6__i5__net25 n7__i5__i6__i5__net25 100.8e-3
rk3911 n8__i5__i6__i5__net25 n9__i5__i6__i5__net25 15.5
rk3912 n6__i5__i6__i5__net21 n9__i5__i6__i5__net21 4.9e-3
rk3913 n8__i5__i6__i5__net21 n9__i5__i6__i5__net21 37.5
rk3914 n9__i5__i8__i10__net25 n7__i5__i8__i10__net25 100.8e-3
rk3915 n8__i5__i8__i10__net25 n9__i5__i8__i10__net25 15.5
rk3916 n6__i5__i8__i10__net21 n9__i5__i8__i10__net21 4.9e-3
rk3917 n8__i5__i8__i10__net21 n9__i5__i8__i10__net21 37.5
rk3919 n1336__vddio n1352__vddio 30.13e-3
rk3920 n1352__vddio n1339__vddio 335.6e-3
rk3921 n1339__vddio n1340__vddio 343.1e-3
rk3922 n1340__vddio n1353__vddio 42.68e-3
rk3923 n1353__vddio n1343__vddio 321.2e-3
rk3924 n1343__vddio n1344__vddio 362.5e-3
rk3925 n1344__vddio n1354__vddio 40.17e-3
rk3926 n1354__vddio n1347__vddio 323.7e-3
rk3927 n1347__vddio n1348__vddio 343.1e-3
rk3928 n1348__vddio n1355__vddio 52.73e-3
rk3929 n1355__vddio n1356__vddio 394.2e-3
rk3930 n1351__vddio n1352__vddio 3.1
rk3931 n1351__vddio n1353__vddio 3.1
rk3932 n1351__vddio n1354__vddio 3.1
rk3933 n1351__vddio n1355__vddio 3.1
rk3934 n803__vss n801__vss 55.24e-3
rk3935 n801__vss n798__vss 365.7e-3
rk3936 n798__vss n804__vss 298.6e-3
rk3937 n804__vss n797__vss 42.68e-3
rk3938 n797__vss n794__vss 365.7e-3
rk3939 n794__vss n805__vss 187.7e-3
rk3940 n805__vss n806__vss 264.6e-3
rk3941 n802__vss n803__vss 3.75
rk3942 n802__vss n804__vss 3.75
rk3943 n802__vss n805__vss 5.7692
rk3946 n2__i5__i6__i5__net24 n3__i5__i6__i5__net24 323.3e-3
rk3947 i5__i6__i5__net24 n2__i5__i6__i5__net24 15.5
rk3948 i5__i6__i5__net23 n2__i5__i6__i5__net23 37.7516
rk3949 n2__i5__i8__i10__net24 n3__i5__i8__i10__net24 323.3e-3
rk3950 i5__i8__i10__net24 n2__i5__i8__i10__net24 15.5
rk3951 i5__i8__i10__net23 n2__i5__i8__i10__net23 37.7516
rk3953 n1075__i1__i14__net1 n1092__i1__i14__net1 210.4e-3
rk3954 n1092__i1__i14__net1 n1076__i1__i14__net1 155.3e-3
rk3955 n1076__i1__i14__net1 n1079__i1__i14__net1 343.1e-3
rk3956 n1079__i1__i14__net1 n1093__i1__i14__net1 226.6e-3
rk3957 n1093__i1__i14__net1 n1080__i1__i14__net1 139.1e-3
rk3958 n1080__i1__i14__net1 n1083__i1__i14__net1 362.5e-3
rk3959 n1083__i1__i14__net1 n1094__i1__i14__net1 223.4e-3
rk3960 n1094__i1__i14__net1 n1084__i1__i14__net1 142.4e-3
rk3961 n1084__i1__i14__net1 n1087__i1__i14__net1 343.1e-3
rk3962 n1087__i1__i14__net1 n1095__i1__i14__net1 239.6e-3
rk3963 n1095__i1__i14__net1 n1088__i1__i14__net1 126.2e-3
rk3965 n1091__i1__i14__net1 n1092__i1__i14__net1 3.1
rk3966 n1091__i1__i14__net1 n1093__i1__i14__net1 3.1
rk3967 n1091__i1__i14__net1 n1094__i1__i14__net1 3.1
rk3968 n1091__i1__i14__net1 n1095__i1__i14__net1 3.1
rk3970 n1099__i1__i14__net1 n1064__i1__i14__net1 12.55e-3
rk3971 n1064__i1__i14__net1 n1067__i1__i14__net1 365.7e-3
rk3972 n1067__i1__i14__net1 n1100__i1__i14__net1 226.6e-3
rk3973 n1100__i1__i14__net1 n1068__i1__i14__net1 116.5e-3
rk3974 n1068__i1__i14__net1 n1071__i1__i14__net1 365.7e-3
rk3975 n1071__i1__i14__net1 n1101__i1__i14__net1 242.8e-3
rk3976 n1101__i1__i14__net1 n1072__i1__i14__net1 119.7e-3
rk3978 n1098__i1__i14__net1 n1099__i1__i14__net1 5.7692
rk3979 n1098__i1__i14__net1 n1100__i1__i14__net1 3.75
rk3980 n1098__i1__i14__net1 n1101__i1__i14__net1 3.75
rk3981 n8__i5__i6__i5__net22 n9__i5__i6__i5__net22 15.9814
rk3982 n9__i5__i6__i5__net22 n10__i5__i6__i5__net22 37.8249
rk3983 n9__i5__i6__i5__net22 n3__i5__i6__i5__net22 22.9156
rk3984 n66__i1__net2 n169__i1__net2 125e-3
rk3985 n68__i1__net2 n170__i1__net2 125e-3
rk3986 n8__i5__i8__i10__net22 n9__i5__i8__i10__net22 15.9814
rk3987 n9__i5__i8__i10__net22 n10__i5__i8__i10__net22 37.8249
rk3988 n9__i5__i8__i10__net22 n3__i5__i8__i10__net22 22.9156
rk3989 n5__i5__i6__i5__net24 n6__i5__i6__i5__net24 350.8e-3
rk3990 n4__i5__i6__i5__net24 n5__i5__i6__i5__net24 15.5
rk3991 n3__i5__i6__i5__net23 n5__i5__i6__i5__net23 4.9e-3
rk3992 n4__i5__i6__i5__net23 n5__i5__i6__i5__net23 37.5
rk3994 n1358__vddio n1360__vddio 30.13e-3
rk3995 n1360__vddio n1361__vddio 335.6e-3
rk3996 n1361__vddio n1362__vddio 343.1e-3
rk3997 n1362__vddio n1363__vddio 42.68e-3
rk3998 n1363__vddio n1364__vddio 321.2e-3
rk3999 n1364__vddio n1365__vddio 362.5e-3
rk4000 n1365__vddio n1366__vddio 40.17e-3
rk4001 n1366__vddio n1367__vddio 323.7e-3
rk4002 n1367__vddio n1368__vddio 343.1e-3
rk4003 n1368__vddio n1369__vddio 52.73e-3
rk4004 n1369__vddio n1370__vddio 394.2e-3
rk4005 n1359__vddio n1360__vddio 3.1
rk4006 n1359__vddio n1363__vddio 3.1
rk4007 n1359__vddio n1366__vddio 3.1
rk4008 n1359__vddio n1369__vddio 3.1
rk4009 n808__vss n809__vss 55.24e-3
rk4010 n809__vss n810__vss 365.7e-3
rk4011 n810__vss n811__vss 298.6e-3
rk4012 n811__vss n812__vss 42.68e-3
rk4013 n812__vss n813__vss 365.7e-3
rk4014 n813__vss n814__vss 187.7e-3
rk4015 n814__vss n815__vss 264.6e-3
rk4016 n807__vss n808__vss 3.75
rk4017 n807__vss n811__vss 3.75
rk4018 n807__vss n814__vss 5.7692
rk4019 n5__i5__i8__i10__net24 n6__i5__i8__i10__net24 350.8e-3
rk4020 n4__i5__i8__i10__net24 n5__i5__i8__i10__net24 15.5
rk4021 n3__i5__i8__i10__net23 n5__i5__i8__i10__net23 4.9e-3
rk4022 n4__i5__i8__i10__net23 n5__i5__i8__i10__net23 37.5
rk4023 n40__i5__i6__net31 n44__i5__i6__net31 500e-3
rk4024 n62__i5__clk_buf n67__i5__clk_buf 500e-3
rk4025 n17__i5__i8__net1 n27__i5__i8__net1 500e-3
rk4026 n15__i5__i8__net2 n35__i5__i8__net2 500e-3
rk4027 n74__i1__net2 n171__i1__net2 125e-3
rk4028 n76__i1__net2 n172__i1__net2 125e-3
rk4030 n1105__i1__i14__net1 n1106__i1__i14__net1 12.55e-3
rk4031 n1106__i1__i14__net1 n1107__i1__i14__net1 365.7e-3
rk4032 n1107__i1__i14__net1 n1108__i1__i14__net1 226.6e-3
rk4033 n1108__i1__i14__net1 n1109__i1__i14__net1 116.5e-3
rk4034 n1109__i1__i14__net1 n1110__i1__i14__net1 365.7e-3
rk4035 n1110__i1__i14__net1 n1111__i1__i14__net1 242.8e-3
rk4036 n1111__i1__i14__net1 n1112__i1__i14__net1 119.7e-3
rk4038 n1104__i1__i14__net1 n1105__i1__i14__net1 5.7692
rk4039 n1104__i1__i14__net1 n1108__i1__i14__net1 3.75
rk4040 n1104__i1__i14__net1 n1111__i1__i14__net1 3.75
rk4042 n1115__i1__i14__net1 n1117__i1__i14__net1 210.4e-3
rk4043 n1117__i1__i14__net1 n1118__i1__i14__net1 155.3e-3
rk4044 n1118__i1__i14__net1 n1119__i1__i14__net1 343.1e-3
rk4045 n1119__i1__i14__net1 n1120__i1__i14__net1 226.6e-3
rk4046 n1120__i1__i14__net1 n1121__i1__i14__net1 139.1e-3
rk4047 n1121__i1__i14__net1 n1122__i1__i14__net1 362.5e-3
rk4048 n1122__i1__i14__net1 n1123__i1__i14__net1 223.4e-3
rk4049 n1123__i1__i14__net1 n1124__i1__i14__net1 142.4e-3
rk4050 n1124__i1__i14__net1 n1125__i1__i14__net1 343.1e-3
rk4051 n1125__i1__i14__net1 n1126__i1__i14__net1 239.6e-3
rk4052 n1126__i1__i14__net1 n1127__i1__i14__net1 126.2e-3
rk4054 n1116__i1__i14__net1 n1117__i1__i14__net1 3.1
rk4055 n1116__i1__i14__net1 n1120__i1__i14__net1 3.1
rk4056 n1116__i1__i14__net1 n1123__i1__i14__net1 3.1
rk4057 n1116__i1__i14__net1 n1126__i1__i14__net1 3.1
rk4058 n9__i5__i6__i5__net24 n7__i5__i6__i5__net24 100.8e-3
rk4059 n8__i5__i6__i5__net24 n9__i5__i6__i5__net24 15.5
rk4060 n6__i5__i6__i5__net23 n9__i5__i6__i5__net23 4.9e-3
rk4061 n8__i5__i6__i5__net23 n9__i5__i6__i5__net23 37.5
rk4062 n8__i5__i8__i10__net24 n9__i5__i8__i10__net24 350.8e-3
rk4063 n7__i5__i8__i10__net24 n8__i5__i8__i10__net24 15.5
rk4064 n6__i5__i8__i10__net23 n8__i5__i8__i10__net23 4.9e-3
rk4065 n7__i5__i8__i10__net23 n8__i5__i8__i10__net23 37.5
rk4066 n86__i1__net2 n177__i1__net2 125e-3
rk4067 n88__i1__net2 n178__i1__net2 125e-3
rk4068 n58__reset n68__reset 250e-3
rk4069 n62__reset n69__reset 250e-3
rk4070 n821__vss n822__vss 55.24e-3
rk4071 n822__vss n823__vss 365.7e-3
rk4072 n823__vss n824__vss 298.6e-3
rk4073 n824__vss n825__vss 42.68e-3
rk4074 n825__vss n826__vss 365.7e-3
rk4075 n826__vss n827__vss 187.7e-3
rk4076 n827__vss n828__vss 264.6e-3
rk4077 n820__vss n821__vss 3.75
rk4078 n820__vss n824__vss 3.75
rk4079 n820__vss n827__vss 5.7692
rk4081 n1379__vddio n1381__vddio 30.13e-3
rk4082 n1381__vddio n1382__vddio 335.6e-3
rk4083 n1382__vddio n1383__vddio 343.1e-3
rk4084 n1383__vddio n1384__vddio 42.68e-3
rk4085 n1384__vddio n1385__vddio 321.2e-3
rk4086 n1385__vddio n1386__vddio 362.5e-3
rk4087 n1386__vddio n1387__vddio 40.17e-3
rk4088 n1387__vddio n1388__vddio 323.7e-3
rk4089 n1388__vddio n1389__vddio 343.1e-3
rk4090 n1389__vddio n1390__vddio 52.73e-3
rk4091 n1390__vddio n1391__vddio 394.2e-3
rk4092 n1380__vddio n1381__vddio 3.1
rk4093 n1380__vddio n1384__vddio 3.1
rk4094 n1380__vddio n1387__vddio 3.1
rk4095 n1380__vddio n1390__vddio 3.1
rk4099 n1144__i1__i14__net1 n1145__i1__i14__net1 12.55e-3
rk4100 n1145__i1__i14__net1 n1146__i1__i14__net1 365.7e-3
rk4101 n1146__i1__i14__net1 n1147__i1__i14__net1 226.6e-3
rk4102 n1147__i1__i14__net1 n1148__i1__i14__net1 116.5e-3
rk4103 n1148__i1__i14__net1 n1149__i1__i14__net1 365.7e-3
rk4104 n1149__i1__i14__net1 n1150__i1__i14__net1 242.8e-3
rk4105 n1150__i1__i14__net1 n1151__i1__i14__net1 119.7e-3
rk4107 n1143__i1__i14__net1 n1144__i1__i14__net1 5.7692
rk4108 n1143__i1__i14__net1 n1147__i1__i14__net1 3.75
rk4109 n1143__i1__i14__net1 n1150__i1__i14__net1 3.75
rk4111 n1154__i1__i14__net1 n1156__i1__i14__net1 210.4e-3
rk4112 n1156__i1__i14__net1 n1157__i1__i14__net1 155.3e-3
rk4113 n1157__i1__i14__net1 n1158__i1__i14__net1 343.1e-3
rk4114 n1158__i1__i14__net1 n1159__i1__i14__net1 226.6e-3
rk4115 n1159__i1__i14__net1 n1160__i1__i14__net1 139.1e-3
rk4116 n1160__i1__i14__net1 n1161__i1__i14__net1 362.5e-3
rk4117 n1161__i1__i14__net1 n1162__i1__i14__net1 223.4e-3
rk4118 n1162__i1__i14__net1 n1163__i1__i14__net1 142.4e-3
rk4119 n1163__i1__i14__net1 n1164__i1__i14__net1 343.1e-3
rk4120 n1164__i1__i14__net1 n1165__i1__i14__net1 239.6e-3
rk4121 n1165__i1__i14__net1 n1166__i1__i14__net1 126.2e-3
rk4123 n1155__i1__i14__net1 n1156__i1__i14__net1 3.1
rk4124 n1155__i1__i14__net1 n1159__i1__i14__net1 3.1
rk4125 n1155__i1__i14__net1 n1162__i1__i14__net1 3.1
rk4126 n1155__i1__i14__net1 n1165__i1__i14__net1 3.1
rk4127 n102__i1__net2 n189__i1__net2 125e-3
rk4128 n104__i1__net2 n190__i1__net2 125e-3
rk4129 n834__vss n835__vss 55.24e-3
rk4130 n835__vss n836__vss 365.7e-3
rk4131 n836__vss n837__vss 298.6e-3
rk4132 n837__vss n838__vss 42.68e-3
rk4133 n838__vss n839__vss 365.7e-3
rk4134 n839__vss n840__vss 187.7e-3
rk4135 n840__vss n841__vss 264.6e-3
rk4136 n833__vss n834__vss 3.75
rk4137 n833__vss n837__vss 3.75
rk4138 n833__vss n840__vss 5.7692
rk4140 n1410__vddio n1412__vddio 30.13e-3
rk4141 n1412__vddio n1413__vddio 335.6e-3
rk4142 n1413__vddio n1414__vddio 343.1e-3
rk4143 n1414__vddio n1415__vddio 42.68e-3
rk4144 n1415__vddio n1416__vddio 321.2e-3
rk4145 n1416__vddio n1417__vddio 362.5e-3
rk4146 n1417__vddio n1418__vddio 40.17e-3
rk4147 n1418__vddio n1419__vddio 323.7e-3
rk4148 n1419__vddio n1420__vddio 343.1e-3
rk4149 n1420__vddio n1421__vddio 52.73e-3
rk4150 n1421__vddio n1422__vddio 394.2e-3
rk4151 n1411__vddio n1412__vddio 3.1
rk4152 n1411__vddio n1415__vddio 3.1
rk4153 n1411__vddio n1418__vddio 3.1
rk4154 n1411__vddio n1421__vddio 3.1
rk4155 n106__i1__net2 n193__i1__net2 125e-3
rk4156 n108__i1__net2 n194__i1__net2 125e-3
rk4157 n4__bufin n5__bufin 18.9833
rk4158 n5__bufin n6__bufin 325.5e-3
rk4159 n6__bufin n7__bufin 420.4e-3
rk4160 n7__bufin n8__bufin 37.828
rk4161 n5__bufin n2__bufin 22.6557
rk4162 n6__bufin n9__bufin 19.0309
rk4163 n7__bufin n10__bufin 15.8422
rk4165 n1182__i1__i14__net1 n1184__i1__i14__net1 210.4e-3
rk4166 n1184__i1__i14__net1 n1185__i1__i14__net1 155.3e-3
rk4167 n1185__i1__i14__net1 n1186__i1__i14__net1 343.1e-3
rk4168 n1186__i1__i14__net1 n1187__i1__i14__net1 226.6e-3
rk4169 n1187__i1__i14__net1 n1188__i1__i14__net1 139.1e-3
rk4170 n1188__i1__i14__net1 n1189__i1__i14__net1 362.5e-3
rk4171 n1189__i1__i14__net1 n1190__i1__i14__net1 223.4e-3
rk4172 n1190__i1__i14__net1 n1191__i1__i14__net1 142.4e-3
rk4173 n1191__i1__i14__net1 n1192__i1__i14__net1 343.1e-3
rk4174 n1192__i1__i14__net1 n1193__i1__i14__net1 239.6e-3
rk4175 n1193__i1__i14__net1 n1194__i1__i14__net1 126.2e-3
rk4177 n1183__i1__i14__net1 n1184__i1__i14__net1 3.1
rk4178 n1183__i1__i14__net1 n1187__i1__i14__net1 3.1
rk4179 n1183__i1__i14__net1 n1190__i1__i14__net1 3.1
rk4180 n1183__i1__i14__net1 n1193__i1__i14__net1 3.1
rk4182 n1198__i1__i14__net1 n1199__i1__i14__net1 12.55e-3
rk4183 n1199__i1__i14__net1 n1200__i1__i14__net1 365.7e-3
rk4184 n1200__i1__i14__net1 n1201__i1__i14__net1 226.6e-3
rk4185 n1201__i1__i14__net1 n1202__i1__i14__net1 116.5e-3
rk4186 n1202__i1__i14__net1 n1203__i1__i14__net1 365.7e-3
rk4187 n1203__i1__i14__net1 n1204__i1__i14__net1 242.8e-3
rk4188 n1204__i1__i14__net1 n1205__i1__i14__net1 119.7e-3
rk4190 n1197__i1__i14__net1 n1198__i1__i14__net1 5.7692
rk4191 n1197__i1__i14__net1 n1201__i1__i14__net1 3.75
rk4192 n1197__i1__i14__net1 n1204__i1__i14__net1 3.75
rk4193 n79__i5__clk4 n89__i5__clk4 22.7255
rk4194 n89__i5__clk4 n90__i5__clk4 184.4e-3
rk4195 n90__i5__clk4 n91__i5__clk4 299.7e-3
rk4196 n91__i5__clk4 n92__i5__clk4 303.9e-3
rk4197 n92__i5__clk4 n93__i5__clk4 37.813
rk4198 n89__i5__clk4 n94__i5__clk4 301.9e-3
rk4199 n90__i5__clk4 n95__i5__clk4 19.0497
rk4200 n91__i5__clk4 n96__i5__clk4 19.0047
rk4201 n92__i5__clk4 n97__i5__clk4 15.8698
rk4202 n114__i1__net2 n197__i1__net2 125e-3
rk4203 n116__i1__net2 n198__i1__net2 125e-3
rk4205 n1431__vddio n1433__vddio 30.13e-3
rk4206 n1433__vddio n1434__vddio 335.6e-3
rk4207 n1434__vddio n1435__vddio 343.1e-3
rk4208 n1435__vddio n1436__vddio 42.68e-3
rk4209 n1436__vddio n1437__vddio 321.2e-3
rk4210 n1437__vddio n1438__vddio 362.5e-3
rk4211 n1438__vddio n1439__vddio 40.17e-3
rk4212 n1439__vddio n1440__vddio 323.7e-3
rk4213 n1440__vddio n1441__vddio 343.1e-3
rk4214 n1441__vddio n1442__vddio 52.73e-3
rk4215 n1442__vddio n1443__vddio 394.2e-3
rk4216 n1432__vddio n1433__vddio 3.1
rk4217 n1432__vddio n1436__vddio 3.1
rk4218 n1432__vddio n1439__vddio 3.1
rk4219 n1432__vddio n1442__vddio 3.1
rk4220 n847__vss n848__vss 55.24e-3
rk4221 n848__vss n849__vss 365.7e-3
rk4222 n849__vss n850__vss 298.6e-3
rk4223 n850__vss n851__vss 42.68e-3
rk4224 n851__vss n852__vss 365.7e-3
rk4225 n852__vss n853__vss 187.7e-3
rk4226 n853__vss n854__vss 264.6e-3
rk4227 n846__vss n847__vss 3.75
rk4228 n846__vss n850__vss 3.75
rk4229 n846__vss n853__vss 5.7692
rk4230 n7__i4__net1 n8__i4__net1 15.8729
rk4231 n8__i4__net1 n9__i4__net1 37.7743
rk4232 n8__i4__net1 n4__i4__net1 45.3022
rk4233 n122__i1__net2 n201__i1__net2 125e-3
rk4234 n124__i1__net2 n202__i1__net2 125e-3
rk4235 n13__i5__i8__net5 n11__i5__i8__net5 31.202
rk4236 n11__i5__i8__net5 n14__i5__i8__net5 42.62e-3
rk4237 n14__i5__i8__net5 n15__i5__i8__net5 279.3e-3
rk4238 n15__i5__i8__net5 n16__i5__i8__net5 75.2422
rk4239 n14__i5__i8__net5 n17__i5__i8__net5 75.2143
rk4240 n15__i5__i8__net5 n18__i5__i8__net5 31.3077
rk4242 n1221__i1__i14__net1 n1223__i1__i14__net1 210.4e-3
rk4243 n1223__i1__i14__net1 n1224__i1__i14__net1 155.3e-3
rk4244 n1224__i1__i14__net1 n1225__i1__i14__net1 343.1e-3
rk4245 n1225__i1__i14__net1 n1226__i1__i14__net1 226.6e-3
rk4246 n1226__i1__i14__net1 n1227__i1__i14__net1 139.1e-3
rk4247 n1227__i1__i14__net1 n1228__i1__i14__net1 362.5e-3
rk4248 n1228__i1__i14__net1 n1229__i1__i14__net1 223.4e-3
rk4249 n1229__i1__i14__net1 n1230__i1__i14__net1 142.4e-3
rk4250 n1230__i1__i14__net1 n1231__i1__i14__net1 343.1e-3
rk4251 n1231__i1__i14__net1 n1232__i1__i14__net1 239.6e-3
rk4252 n1232__i1__i14__net1 n1233__i1__i14__net1 126.2e-3
rk4254 n1222__i1__i14__net1 n1223__i1__i14__net1 3.1
rk4255 n1222__i1__i14__net1 n1226__i1__i14__net1 3.1
rk4256 n1222__i1__i14__net1 n1229__i1__i14__net1 3.1
rk4257 n1222__i1__i14__net1 n1232__i1__i14__net1 3.1
rk4259 n1237__i1__i14__net1 n1238__i1__i14__net1 12.55e-3
rk4260 n1238__i1__i14__net1 n1239__i1__i14__net1 365.7e-3
rk4261 n1239__i1__i14__net1 n1240__i1__i14__net1 226.6e-3
rk4262 n1240__i1__i14__net1 n1241__i1__i14__net1 116.5e-3
rk4263 n1241__i1__i14__net1 n1242__i1__i14__net1 365.7e-3
rk4264 n1242__i1__i14__net1 n1243__i1__i14__net1 242.8e-3
rk4265 n1243__i1__i14__net1 n1244__i1__i14__net1 119.7e-3
rk4267 n1236__i1__i14__net1 n1237__i1__i14__net1 5.7692
rk4268 n1236__i1__i14__net1 n1240__i1__i14__net1 3.75
rk4269 n1236__i1__i14__net1 n1243__i1__i14__net1 3.75
rk4270 n134__i1__net2 n205__i1__net2 125e-3
rk4271 n136__i1__net2 n206__i1__net2 125e-3
rk4273 n1452__vddio n1454__vddio 30.13e-3
rk4274 n1454__vddio n1455__vddio 335.6e-3
rk4275 n1455__vddio n1456__vddio 343.1e-3
rk4276 n1456__vddio n1457__vddio 42.68e-3
rk4277 n1457__vddio n1458__vddio 321.2e-3
rk4278 n1458__vddio n1459__vddio 362.5e-3
rk4279 n1459__vddio n1460__vddio 40.17e-3
rk4280 n1460__vddio n1461__vddio 323.7e-3
rk4281 n1461__vddio n1462__vddio 343.1e-3
rk4282 n1462__vddio n1463__vddio 52.73e-3
rk4283 n1463__vddio n1464__vddio 394.2e-3
rk4284 n1453__vddio n1454__vddio 3.1
rk4285 n1453__vddio n1457__vddio 3.1
rk4286 n1453__vddio n1460__vddio 3.1
rk4287 n1453__vddio n1463__vddio 3.1
rk4288 n860__vss n861__vss 55.24e-3
rk4289 n861__vss n862__vss 365.7e-3
rk4290 n862__vss n863__vss 298.6e-3
rk4291 n863__vss n864__vss 42.68e-3
rk4292 n864__vss n865__vss 365.7e-3
rk4293 n865__vss n866__vss 187.7e-3
rk4294 n866__vss n867__vss 264.6e-3
rk4295 n859__vss n860__vss 3.75
rk4296 n859__vss n863__vss 3.75
rk4297 n859__vss n866__vss 5.7692
rk4298 n87__i5__clk4 n101__i5__clk4 500e-3
rk4299 n14__piso_out n15__piso_out 15.9076
rk4300 n15__piso_out n6__piso_out 185e-3
rk4302 n15__piso_out n17__piso_out 37.7974
rk4303 n138__i1__net2 n209__i1__net2 125e-3
rk4304 n140__i1__net2 n210__i1__net2 125e-3
rk4305 n32__i5__i8__net2 n37__i5__i8__net2 502.5e-3
rk4307 n1261__i1__i14__net1 n1262__i1__i14__net1 12.55e-3
rk4308 n1262__i1__i14__net1 n1263__i1__i14__net1 365.7e-3
rk4309 n1263__i1__i14__net1 n1264__i1__i14__net1 226.6e-3
rk4310 n1264__i1__i14__net1 n1265__i1__i14__net1 116.5e-3
rk4311 n1265__i1__i14__net1 n1266__i1__i14__net1 365.7e-3
rk4312 n1266__i1__i14__net1 n1267__i1__i14__net1 242.8e-3
rk4313 n1267__i1__i14__net1 n1268__i1__i14__net1 119.7e-3
rk4315 n1260__i1__i14__net1 n1261__i1__i14__net1 5.7692
rk4316 n1260__i1__i14__net1 n1264__i1__i14__net1 3.75
rk4317 n1260__i1__i14__net1 n1267__i1__i14__net1 3.75
rk4319 n1271__i1__i14__net1 n1273__i1__i14__net1 210.4e-3
rk4320 n1273__i1__i14__net1 n1274__i1__i14__net1 155.3e-3
rk4321 n1274__i1__i14__net1 n1275__i1__i14__net1 343.1e-3
rk4322 n1275__i1__i14__net1 n1276__i1__i14__net1 226.6e-3
rk4323 n1276__i1__i14__net1 n1277__i1__i14__net1 139.1e-3
rk4324 n1277__i1__i14__net1 n1278__i1__i14__net1 362.5e-3
rk4325 n1278__i1__i14__net1 n1279__i1__i14__net1 223.4e-3
rk4326 n1279__i1__i14__net1 n1280__i1__i14__net1 142.4e-3
rk4327 n1280__i1__i14__net1 n1281__i1__i14__net1 343.1e-3
rk4328 n1281__i1__i14__net1 n1282__i1__i14__net1 239.6e-3
rk4329 n1282__i1__i14__net1 n1283__i1__i14__net1 126.2e-3
rk4331 n1272__i1__i14__net1 n1273__i1__i14__net1 3.1
rk4332 n1272__i1__i14__net1 n1276__i1__i14__net1 3.1
rk4333 n1272__i1__i14__net1 n1279__i1__i14__net1 3.1
rk4334 n1272__i1__i14__net1 n1282__i1__i14__net1 3.1
rk4337 n881__vss n878__vss 55.24e-3
rk4338 n878__vss n877__vss 365.7e-3
rk4339 n877__vss n882__vss 298.6e-3
rk4340 n882__vss n874__vss 42.68e-3
rk4341 n874__vss n873__vss 365.7e-3
rk4342 n873__vss n883__vss 187.7e-3
rk4343 n883__vss n884__vss 264.6e-3
rk4344 n880__vss n881__vss 3.75
rk4345 n880__vss n882__vss 3.75
rk4346 n880__vss n883__vss 5.7692
rk4348 n1473__vddio n1488__vddio 30.13e-3
rk4349 n1488__vddio n1474__vddio 335.6e-3
rk4350 n1474__vddio n1477__vddio 343.1e-3
rk4351 n1477__vddio n1489__vddio 42.68e-3
rk4352 n1489__vddio n1478__vddio 321.2e-3
rk4353 n1478__vddio n1481__vddio 362.5e-3
rk4354 n1481__vddio n1490__vddio 40.17e-3
rk4355 n1490__vddio n1482__vddio 323.7e-3
rk4356 n1482__vddio n1485__vddio 343.1e-3
rk4357 n1485__vddio n1491__vddio 52.73e-3
rk4358 n1491__vddio n1492__vddio 394.2e-3
rk4359 n1487__vddio n1488__vddio 3.1
rk4360 n1487__vddio n1489__vddio 3.1
rk4361 n1487__vddio n1490__vddio 3.1
rk4362 n1487__vddio n1491__vddio 3.1
rk4363 n4__piso_outinv n2__piso_outinv 31.2855
rk4364 n2__piso_outinv n5__piso_outinv 223e-3
rk4365 n5__piso_outinv n6__piso_outinv 75.3031
rk4366 n2__piso_outinv n7__piso_outinv 75.2361
rk4367 n5__piso_outinv n8__piso_outinv 31.3339
rk4368 n154__i1__net2 n217__i1__net2 125e-3
rk4369 n156__i1__net2 n218__i1__net2 125e-3
rk4370 n4__i5__i8__i8__net1 n5__i5__i8__i8__net1 15.8129
rk4371 n5__i5__i8__i8__net1 n6__i5__i8__i8__net1 75.3643
rk4372 n5__i5__i8__i8__net1 n2__i5__i8__i8__net1 45.336
rk4374 n1326__i1__i14__net1 n1298__i1__i14__net1 12.55e-3
rk4375 n1298__i1__i14__net1 n1301__i1__i14__net1 365.7e-3
rk4376 n1301__i1__i14__net1 n1327__i1__i14__net1 226.6e-3
rk4377 n1327__i1__i14__net1 n1302__i1__i14__net1 116.5e-3
rk4378 n1302__i1__i14__net1 n1305__i1__i14__net1 365.7e-3
rk4379 n1305__i1__i14__net1 n1328__i1__i14__net1 242.8e-3
rk4380 n1328__i1__i14__net1 n1306__i1__i14__net1 119.7e-3
rk4382 n1325__i1__i14__net1 n1326__i1__i14__net1 5.7692
rk4383 n1325__i1__i14__net1 n1327__i1__i14__net1 3.75
rk4384 n1325__i1__i14__net1 n1328__i1__i14__net1 3.75
rk4386 n1309__i1__i14__net1 n1332__i1__i14__net1 210.4e-3
rk4387 n1332__i1__i14__net1 n1310__i1__i14__net1 155.3e-3
rk4388 n1310__i1__i14__net1 n1313__i1__i14__net1 343.1e-3
rk4389 n1313__i1__i14__net1 n1333__i1__i14__net1 226.6e-3
rk4390 n1333__i1__i14__net1 n1314__i1__i14__net1 139.1e-3
rk4391 n1314__i1__i14__net1 n1317__i1__i14__net1 362.5e-3
rk4392 n1317__i1__i14__net1 n1334__i1__i14__net1 223.4e-3
rk4393 n1334__i1__i14__net1 n1318__i1__i14__net1 142.4e-3
rk4394 n1318__i1__i14__net1 n1321__i1__i14__net1 343.1e-3
rk4395 n1321__i1__i14__net1 n1335__i1__i14__net1 239.6e-3
rk4396 n1335__i1__i14__net1 n1322__i1__i14__net1 126.2e-3
rk4398 n1331__i1__i14__net1 n1332__i1__i14__net1 3.1
rk4399 n1331__i1__i14__net1 n1333__i1__i14__net1 3.1
rk4400 n1331__i1__i14__net1 n1334__i1__i14__net1 3.1
rk4401 n1331__i1__i14__net1 n1335__i1__i14__net1 3.1
rk4402 n44__shift n45__shift 15.8284
rk4403 n45__shift n46__shift 37.7016
rk4404 n182__i1__net2 n221__i1__net2 125e-3
rk4405 n184__i1__net2 n222__i1__net2 125e-3
rk4406 n909__vss n891__vss 55.24e-3
rk4407 n891__vss n890__vss 365.7e-3
rk4408 n890__vss n910__vss 298.6e-3
rk4409 n910__vss n887__vss 42.68e-3
rk4410 n887__vss n886__vss 365.7e-3
rk4411 n886__vss n911__vss 187.7e-3
rk4412 n911__vss n893__vss 264.6e-3
rk4413 n908__vss n909__vss 3.75
rk4414 n908__vss n910__vss 3.75
rk4415 n908__vss n911__vss 5.7692
rk4417 n1494__vddio n1524__vddio 30.13e-3
rk4418 n1524__vddio n1495__vddio 335.6e-3
rk4419 n1495__vddio n1498__vddio 343.1e-3
rk4420 n1498__vddio n1525__vddio 42.68e-3
rk4421 n1525__vddio n1499__vddio 321.2e-3
rk4422 n1499__vddio n1502__vddio 362.5e-3
rk4423 n1502__vddio n1526__vddio 40.17e-3
rk4424 n1526__vddio n1503__vddio 323.7e-3
rk4425 n1503__vddio n1506__vddio 343.1e-3
rk4426 n1506__vddio n1527__vddio 52.73e-3
rk4427 n1527__vddio n1507__vddio 394.2e-3
rk4428 n1523__vddio n1524__vddio 3.1
rk4429 n1523__vddio n1525__vddio 3.1
rk4430 n1523__vddio n1526__vddio 3.1
rk4431 n1523__vddio n1527__vddio 3.1
rk4432 n181__vdd n183__vdd 16.0582
rk4433 n183__vdd n184__vdd 92.15e-3
rk4434 n184__vdd n185__vdd 100.2e-3
rk4435 n185__vdd n186__vdd 8.034e-3
rk4436 n186__vdd n187__vdd 43.22e-3
rk4437 n187__vdd n188__vdd 73.73e-3
rk4438 n188__vdd n189__vdd 246.6e-3
rk4439 n189__vdd n190__vdd 127e-3
rk4440 n190__vdd n191__vdd 124.5e-3
rk4441 n191__vdd n192__vdd 106.8e-3
rk4442 n192__vdd n193__vdd 8.034e-3
rk4443 n193__vdd n194__vdd 95.88e-3
rk4444 n194__vdd n195__vdd 138.2e-3
rk4445 n195__vdd n196__vdd 169e-3
rk4446 n196__vdd n197__vdd 16.85e-3
rk4447 n197__vdd n198__vdd 92.77e-3
rk4448 n198__vdd n199__vdd 31.69e-3
rk4449 n199__vdd n200__vdd 105.3e-3
rk4450 n200__vdd n201__vdd 8.034e-3
rk4451 n201__vdd n202__vdd 43.22e-3
rk4452 n202__vdd n160__vdd 72.24e-3
rk4453 n160__vdd n158__vdd 43.72e-3
rk4454 n158__vdd n154__vdd 44.31e-3
rk4456 n154__vdd n204__vdd 6.171e-3
rk4457 n204__vdd n205__vdd 45.39e-3
rk4458 n205__vdd n206__vdd 50.31e-3
rk4459 n206__vdd n207__vdd 110.9e-3
rk4460 n207__vdd n208__vdd 21.26e-3
rk4461 n208__vdd n209__vdd 207.2e-3
rk4462 n209__vdd n210__vdd 191.8e-3
rk4463 n210__vdd n211__vdd 163.1e-3
rk4464 n211__vdd n212__vdd 221.1e-3
rk4465 n212__vdd n213__vdd 10.76e-3
rk4466 n213__vdd n214__vdd 75.06e-3
rk4467 n214__vdd n215__vdd 54.18e-3
rk4468 n215__vdd n216__vdd 171.4e-3
rk4469 n216__vdd n217__vdd 168.9e-3
rk4470 n217__vdd n218__vdd 15.03e-3
rk4471 n218__vdd n219__vdd 127.4e-3
rk4472 n219__vdd n220__vdd 10.69e-3
rk4473 n220__vdd n222__vdd 166.5e-3
rk4474 n222__vdd n223__vdd 19.5e-3
rk4475 n223__vdd n224__vdd 147.1e-3
rk4476 n224__vdd n225__vdd 140.6e-3
rk4477 n225__vdd n226__vdd 10.58e-3
rk4478 n226__vdd n227__vdd 34.09e-3
rk4479 n227__vdd n229__vdd 134.4e-3
rk4480 n229__vdd n230__vdd 132e-3
rk4481 n230__vdd n231__vdd 11.07e-3
rk4482 n231__vdd n232__vdd 72.07e-3
rk4483 n232__vdd n234__vdd 106.8e-3
rk4484 n234__vdd n235__vdd 132e-3
rk4485 n235__vdd n236__vdd 11.07e-3
rk4486 n236__vdd n238__vdd 85.8e-3
rk4487 n238__vdd n239__vdd 13.7e-3
rk4488 n239__vdd n240__vdd 150.7e-3
rk4489 n240__vdd n241__vdd 138.8e-3
rk4490 n241__vdd n242__vdd 59.09e-3
rk4491 n242__vdd n243__vdd 11.21e-3
rk4492 n243__vdd n244__vdd 164.4e-3
rk4493 n244__vdd n245__vdd 138.8e-3
rk4494 n245__vdd n246__vdd 34.18e-3
rk4495 n246__vdd n247__vdd 32.38e-3
rk4496 n247__vdd n248__vdd 164.4e-3
rk4497 n248__vdd n249__vdd 151.9e-3
rk4498 n249__vdd n250__vdd 57.28e-3
rk4499 n250__vdd n251__vdd 164.4e-3
rk4500 n251__vdd n252__vdd 127e-3
rk4501 n252__vdd n253__vdd 77.83e-3
rk4502 n253__vdd n254__vdd 11.05e-3
rk4503 n254__vdd n255__vdd 2.5894
rk4504 n255__vdd n257__vdd 45.32e-3
rk4505 n257__vdd n258__vdd 271.5e-3
rk4506 n258__vdd n259__vdd 571.4e-3
rk4507 n259__vdd n260__vdd 688.1e-3
rk4508 n260__vdd n261__vdd 293.6e-3
rk4509 n261__vdd n262__vdd 572.9e-3
rk4510 n262__vdd n263__vdd 688.1e-3
rk4511 n263__vdd n264__vdd 278.2e-3
rk4512 n264__vdd n265__vdd 572.9e-3
rk4513 n265__vdd n266__vdd 688.1e-3
rk4514 n266__vdd n267__vdd 293.6e-3
rk4515 n267__vdd n268__vdd 572.9e-3
rk4516 n183__vdd n269__vdd 15.9963
rk4517 n185__vdd n270__vdd 31.508
rk4518 n187__vdd n271__vdd 31.4959
rk4519 n190__vdd n272__vdd 15.9932
rk4520 n191__vdd n273__vdd 15.9698
rk4521 n192__vdd n274__vdd 31.508
rk4522 n195__vdd n275__vdd 31.5104
rk4523 n196__vdd n276__vdd 15.9604
rk4524 n199__vdd n277__vdd 15.9698
rk4525 n200__vdd n278__vdd 31.508
rk4526 n202__vdd n279__vdd 31.4959
rk4527 n205__vdd n280__vdd 15.9365
rk4528 n206__vdd n281__vdd 15.9381
rk4529 n208__vdd n282__vdd 31.2407
rk4530 n209__vdd n283__vdd 31.1765
rk4531 n211__vdd n284__vdd 31.1765
rk4532 n213__vdd n285__vdd 31.2557
rk4533 n216__vdd n286__vdd 31.3361
rk4534 n220__vdd n287__vdd 31.253
rk4535 n226__vdd n288__vdd 31.2564
rk4536 n231__vdd n289__vdd 31.2522
rk4537 n236__vdd n290__vdd 31.2522
rk4538 n240__vdd n291__vdd 31.3865
rk4539 n241__vdd n292__vdd 31.4138
rk4540 n244__vdd n293__vdd 31.3865
rk4541 n245__vdd n294__vdd 31.4138
rk4542 n248__vdd n295__vdd 31.3865
rk4543 n249__vdd n296__vdd 31.4524
rk4544 n251__vdd n297__vdd 31.3865
rk4545 n252__vdd n298__vdd 31.4118
rk4546 n254__vdd n299__vdd 31.2551
rk4547 n255__vdd n300__vdd 31.2229
rk4548 n258__vdd n301__vdd 31.3813
rk4549 n259__vdd n302__vdd 31.4122
rk4550 n261__vdd n303__vdd 31.4034
rk4551 n262__vdd n304__vdd 31.4122
rk4552 n264__vdd n305__vdd 31.4034
rk4553 n265__vdd n306__vdd 31.4122
rk4554 n267__vdd n307__vdd 31.4034
rk4555 n268__vdd n308__vdd 31.4122
rk4556 n268__vdd n309__vdd 688.1e-3
rk4557 n309__vdd n310__vdd 361e-3
rk4558 n310__vdd n311__vdd 31.2394
rk4559 n310__vdd n313__vdd 28.25e-3
rk4560 n313__vdd n314__vdd 416.8e-3
rk4561 n314__vdd n315__vdd 669.8e-3
rk4562 n315__vdd n316__vdd 31.2665
rk4563 n315__vdd n318__vdd 35.8e-3
rk4564 n318__vdd n319__vdd 416.8e-3
rk4565 n319__vdd n320__vdd 620.7e-3
rk4566 n320__vdd n321__vdd 31.2135
rk4567 n320__vdd n323__vdd 35.41e-3
rk4568 n323__vdd n324__vdd 466.6e-3
rk4569 n324__vdd n325__vdd 552.9e-3
rk4570 n325__vdd n326__vdd 571.3e-3
rk4571 n326__vdd n327__vdd 31.2135
rk4572 n326__vdd n329__vdd 35.41e-3
rk4573 n329__vdd n330__vdd 466.6e-3
rk4574 n330__vdd n331__vdd 554.4e-3
rk4575 n331__vdd n332__vdd 542.4e-3
rk4576 n332__vdd n333__vdd 31.4623
rk4577 n332__vdd n334__vdd 178e-3
rk4578 n334__vdd n335__vdd 33.12e-3
rk4579 n335__vdd n336__vdd 31.4739
rk4580 n335__vdd n337__vdd 348.8e-3
rk4581 n337__vdd n338__vdd 31.4946
rk4582 n337__vdd n46__vdd 166.7e-3
rk4583 n46__vdd n339__vdd 137.1e-3
rk4584 n339__vdd n340__vdd 660.8e-3
rk4585 n340__vdd n341__vdd 15.9367
rk4586 n340__vdd n342__vdd 499.9e-3
rk4587 n342__vdd n343__vdd 99.78e-3
rk4588 n343__vdd n344__vdd 15.942
rk4589 n343__vdd n345__vdd 650.1e-3
rk4590 n345__vdd n346__vdd 270.1e-3
rk4591 n346__vdd n347__vdd 31.4946
rk4592 n346__vdd n348__vdd 324.8e-3
rk4593 n348__vdd n349__vdd 660.8e-3
rk4594 n349__vdd n350__vdd 15.9367
rk4595 n349__vdd n351__vdd 499.9e-3
rk4596 n351__vdd n352__vdd 99.78e-3
rk4597 n352__vdd n353__vdd 15.942
rk4598 n352__vdd n354__vdd 650.1e-3
rk4599 n354__vdd n355__vdd 277.8e-3
rk4600 n355__vdd n356__vdd 31.4946
rk4601 n355__vdd n357__vdd 324.8e-3
rk4602 n357__vdd n358__vdd 660.8e-3
rk4603 n358__vdd n359__vdd 15.9367
rk4604 n358__vdd n360__vdd 499.9e-3
rk4605 n360__vdd n361__vdd 99.78e-3
rk4606 n361__vdd n362__vdd 15.942
rk4607 n361__vdd n363__vdd 650.1e-3
rk4608 n363__vdd n364__vdd 247.1e-3
rk4609 n364__vdd n365__vdd 15.904
rk4610 n364__vdd n366__vdd 258.6e-3
rk4611 n366__vdd n367__vdd 40.81e-3
rk4612 n367__vdd n368__vdd 15.904
rk4613 n367__vdd n369__vdd 207.2e-3
rk4614 n369__vdd n370__vdd 15.9024
rk4615 n369__vdd n371__vdd 177.8e-3
rk4616 n371__vdd n372__vdd 31.1775
rk4617 n371__vdd n373__vdd 149.5e-3
rk4618 n373__vdd n374__vdd 31.2143
rk4619 n373__vdd n375__vdd 31.3471
rk4620 n182__vdd n183__vdd 7.5
rk4621 n182__vdd n186__vdd 9.375
rk4622 n182__vdd n188__vdd 15
rk4623 n182__vdd n190__vdd 3.75
rk4624 n182__vdd n193__vdd 9.375
rk4625 n182__vdd n195__vdd 15
rk4626 n182__vdd n197__vdd 3.75
rk4627 n182__vdd n201__vdd 9.375
rk4628 n182__vdd n204__vdd 5
rk4629 n182__vdd n207__vdd 25
rk4630 n182__vdd n210__vdd 5.3571
rk4631 n182__vdd n212__vdd 25
rk4632 n47__vdd n214__vdd 12.5e-3
rk4633 n182__vdd n215__vdd 7.5
rk4634 n182__vdd n216__vdd 25
rk4635 n49__vdd n217__vdd 12.5e-3
rk4636 n182__vdd n218__vdd 7.5
rk4637 n182__vdd n219__vdd 25
rk4638 n221__vdd n222__vdd 7.5
rk4639 n51__vdd n223__vdd 12.5e-3
rk4640 n221__vdd n224__vdd 7.5
rk4641 n221__vdd n225__vdd 25
rk4642 n53__vdd n227__vdd 12.5e-3
rk4643 n228__vdd n229__vdd 7.5
rk4644 n228__vdd n230__vdd 25
rk4645 n55__vdd n232__vdd 12.5e-3
rk4646 n233__vdd n234__vdd 7.5
rk4647 n233__vdd n235__vdd 25
rk4648 n237__vdd n238__vdd 37.5
rk4649 n57__vdd n239__vdd 12.5e-3
rk4650 n237__vdd n240__vdd 3.75
rk4651 n59__vdd n242__vdd 12.5e-3
rk4652 n237__vdd n243__vdd 37.5
rk4653 n237__vdd n244__vdd 3.75
rk4654 n61__vdd n246__vdd 12.5e-3
rk4655 n237__vdd n247__vdd 37.5
rk4656 n237__vdd n248__vdd 3.75
rk4657 n63__vdd n249__vdd 12.5e-3
rk4658 n237__vdd n250__vdd 37.5
rk4659 n237__vdd n251__vdd 3.75
rk4660 n65__vdd n252__vdd 12.5e-3
rk4661 n237__vdd n253__vdd 25
rk4662 n256__vdd n257__vdd 25
rk4663 n256__vdd n259__vdd 3.75
rk4664 n256__vdd n260__vdd 37.5
rk4665 n256__vdd n262__vdd 3.75
rk4666 n256__vdd n263__vdd 37.5
rk4667 n256__vdd n265__vdd 3.75
rk4668 n256__vdd n266__vdd 37.5
rk4669 n256__vdd n268__vdd 3.75
rk4670 n256__vdd n309__vdd 37.5
rk4671 n312__vdd n313__vdd 25
rk4672 n312__vdd n314__vdd 7.5
rk4673 n317__vdd n318__vdd 25
rk4674 n317__vdd n319__vdd 7.5
rk4675 n322__vdd n323__vdd 25
rk4676 n322__vdd n324__vdd 7.5
rk4677 n322__vdd n325__vdd 7.5
rk4678 n328__vdd n329__vdd 25
rk4679 n328__vdd n330__vdd 7.5
rk4680 n328__vdd n331__vdd 7.5
rk4681 n328__vdd n334__vdd 9.375
rk4682 n328__vdd n339__vdd 6.25
rk4683 n328__vdd n342__vdd 3.75
rk4684 n328__vdd n345__vdd 15
rk4685 n328__vdd n348__vdd 6.25
rk4686 n328__vdd n351__vdd 3.75
rk4687 n328__vdd n354__vdd 15
rk4688 n328__vdd n357__vdd 6.25
rk4689 n328__vdd n360__vdd 3.75
rk4690 n328__vdd n363__vdd 15
rk4691 n328__vdd n366__vdd 7.5
rk4692 n328__vdd n373__vdd 9.375
rk4693 n1632__vddio n1633__vddio 57.6e-3
rk4694 n1633__vddio n1634__vddio 142.3e-3
rk4695 n1634__vddio n1635__vddio 142.3e-3
rk4696 n1635__vddio n1636__vddio 183e-3
rk4697 n1636__vddio n1637__vddio 196.5e-3
rk4698 n1637__vddio n1638__vddio 128.8e-3
rk4699 n1638__vddio n1639__vddio 250.7e-3
rk4700 n1639__vddio n1640__vddio 74.54e-3
rk4701 n1640__vddio n1641__vddio 304.9e-3
rk4702 n1641__vddio n1642__vddio 20.33e-3
rk4703 n1642__vddio n1643__vddio 325.3e-3
rk4704 n1643__vddio n1644__vddio 33.88e-3
rk4705 n1644__vddio n1645__vddio 291.4e-3
rk4706 n1645__vddio n1646__vddio 88.09e-3
rk4707 n1646__vddio n1647__vddio 237.2e-3
rk4708 n1647__vddio n1648__vddio 142.3e-3
rk4709 n1648__vddio n1649__vddio 183e-3
rk4710 n1649__vddio n1650__vddio 196.5e-3
rk4711 n1650__vddio n1651__vddio 128.8e-3
rk4712 n1651__vddio n1652__vddio 250.7e-3
rk4713 n1652__vddio n1653__vddio 74.54e-3
rk4714 n1653__vddio n1654__vddio 304.9e-3
rk4715 n1654__vddio n1655__vddio 20.33e-3
rk4716 n1655__vddio n1656__vddio 325.3e-3
rk4717 n1656__vddio n1657__vddio 33.88e-3
rk4718 n1657__vddio n1658__vddio 291.4e-3
rk4719 n1658__vddio n1659__vddio 88.09e-3
rk4720 n1659__vddio n1660__vddio 237.2e-3
rk4721 n1660__vddio n1661__vddio 142.3e-3
rk4722 n1661__vddio n1662__vddio 183e-3
rk4723 n1662__vddio n1663__vddio 196.5e-3
rk4724 n1663__vddio n1664__vddio 128.8e-3
rk4725 n1664__vddio n1665__vddio 250.7e-3
rk4726 n1665__vddio n1666__vddio 74.54e-3
rk4727 n1666__vddio n1667__vddio 304.9e-3
rk4728 n1667__vddio n1631__vddio 1.2703
rk4729 n1631__vddio n1632__vddio 5
rk4730 n1529__vddio n1633__vddio 16.67e-3
rk4731 n1631__vddio n1634__vddio 1.25
rk4732 n1533__vddio n1635__vddio 8.333e-3
rk4733 n1631__vddio n1636__vddio 1.25
rk4734 n1538__vddio n1637__vddio 8.333e-3
rk4735 n1631__vddio n1638__vddio 1.25
rk4736 n1543__vddio n1639__vddio 8.333e-3
rk4737 n1631__vddio n1640__vddio 1.25
rk4738 n1547__vddio n1641__vddio 8.333e-3
rk4739 n1631__vddio n1642__vddio 1.25
rk4740 n1631__vddio n1643__vddio 1.25
rk4741 n1551__vddio n1644__vddio 8.333e-3
rk4742 n1631__vddio n1645__vddio 1.25
rk4743 n1555__vddio n1646__vddio 8.333e-3
rk4744 n1631__vddio n1647__vddio 1.25
rk4745 n1559__vddio n1648__vddio 8.333e-3
rk4746 n1631__vddio n1649__vddio 1.25
rk4747 n1563__vddio n1650__vddio 8.333e-3
rk4748 n1631__vddio n1651__vddio 1.25
rk4749 n1567__vddio n1652__vddio 8.333e-3
rk4750 n1631__vddio n1653__vddio 1.25
rk4751 n1571__vddio n1654__vddio 8.333e-3
rk4752 n1631__vddio n1655__vddio 1.25
rk4753 n1631__vddio n1656__vddio 1.25
rk4754 n1575__vddio n1657__vddio 8.333e-3
rk4755 n1631__vddio n1658__vddio 1.25
rk4756 n1579__vddio n1659__vddio 8.333e-3
rk4757 n1631__vddio n1660__vddio 1.25
rk4758 n1583__vddio n1661__vddio 8.333e-3
rk4759 n1631__vddio n1662__vddio 1.25
rk4760 n1587__vddio n1663__vddio 8.333e-3
rk4761 n1631__vddio n1664__vddio 1.25
rk4762 n1591__vddio n1665__vddio 8.333e-3
rk4763 n1631__vddio n1666__vddio 1.25
rk4764 n1595__vddio n1667__vddio 8.333e-3
rk4765 n1014__vss n1015__vss 47.96e-3
rk4766 n1015__vss n1016__vss 150.4e-3
rk4767 n1016__vss n1017__vss 134.2e-3
rk4768 n1017__vss n1018__vss 191.1e-3
rk4769 n1018__vss n1019__vss 59.63e-3
rk4770 n1019__vss n1020__vss 128.8e-3
rk4771 n1020__vss n1021__vss 136.9e-3
rk4772 n1021__vss n1022__vss 177.5e-3
rk4773 n1022__vss n1023__vss 65.05e-3
rk4774 n1023__vss n1024__vss 82.67e-3
rk4775 n1024__vss n1025__vss 257.5e-3
rk4776 n1025__vss n1026__vss 39.3e-3
rk4777 n1026__vss n1027__vss 28.46e-3
rk4778 n1027__vss n1028__vss 110.5e-3
rk4779 n1028__vss n1029__vss 214.8e-3
rk4780 n1029__vss n1030__vss 5.346e-3
rk4781 n1030__vss n1031__vss 299.5e-3
rk4782 n1031__vss n1032__vss 79.96e-3
rk4783 n1032__vss n1033__vss 245.3e-3
rk4784 n1033__vss n1034__vss 61.67e-3
rk4785 n1034__vss n1035__vss 72.51e-3
rk4786 n1035__vss n1036__vss 191.1e-3
rk4787 n1036__vss n1037__vss 188.4e-3
rk4788 n1037__vss n1038__vss 60.31e-3
rk4789 n1038__vss n1039__vss 76.57e-3
rk4790 n1039__vss n1040__vss 242.6e-3
rk4791 n1040__vss n1041__vss 82.67e-3
rk4792 n1041__vss n1042__vss 122.7e-3
rk4793 n1042__vss n1043__vss 174.2e-3
rk4794 n1043__vss n1044__vss 28.46e-3
rk4795 n1044__vss n1045__vss 160.6e-3
rk4796 n1045__vss n1046__vss 164.7e-3
rk4797 n1046__vss n1047__vss 25.75e-3
rk4798 n1047__vss n1048__vss 132.8e-3
rk4799 n1048__vss n1049__vss 166.7e-3
rk4800 n1049__vss n1050__vss 79.96e-3
rk4801 n1050__vss n1051__vss 174.2e-3
rk4802 n1051__vss n1052__vss 71.15e-3
rk4803 n1052__vss n1053__vss 134.2e-3
rk4804 n1053__vss n1054__vss 191.1e-3
rk4805 n1054__vss n1055__vss 188.4e-3
rk4806 n1055__vss n1056__vss 136.9e-3
rk4807 n1056__vss n1057__vss 88.02e-3
rk4808 n1057__vss n1058__vss 154.4e-3
rk4809 n1058__vss n1059__vss 82.67e-3
rk4810 n1059__vss n1060__vss 296.8e-3
rk4811 n1060__vss n1013__vss 1.0618
rk4812 n1057__vss n1061__vss 613.7e-3
rk4813 n1061__vss n1062__vss 184.3e-3
rk4814 n1062__vss n1063__vss 48.49e-3
rk4815 n1063__vss n1064__vss 628.3e-3
rk4816 n1064__vss n1065__vss 672.8e-3
rk4817 n1065__vss n1066__vss 147.4e-3
rk4818 n1066__vss n1067__vss 75.4606
rk4819 n1061__vss n1068__vss 104.7e-3
rk4820 n1068__vss n1069__vss 75.4253
rk4821 n1063__vss n1070__vss 19.1362
rk4822 n1064__vss n1071__vss 75.4386
rk4823 n1065__vss n1072__vss 75.4748
rk4824 n1068__vss n1073__vss 571.3e-3
rk4825 n1073__vss n1074__vss 75.4386
rk4826 n1073__vss n1075__vss 628.3e-3
rk4827 n1075__vss n1076__vss 19.1362
rk4828 n1075__vss n1077__vss 48.49e-3
rk4829 n1077__vss n1078__vss 159.5e-3
rk4830 n1078__vss n1079__vss 290.3e-3
rk4831 n1078__vss n1080__vss 115.8e-3
rk4832 n1080__vss n1081__vss 75.4253
rk4833 n1079__vss n1054__vss 304.8e-3
rk4834 n1080__vss n1082__vss 571.3e-3
rk4835 n1082__vss n1083__vss 75.4386
rk4836 n1082__vss n1084__vss 628.3e-3
rk4837 n1084__vss n1085__vss 19.1362
rk4838 n1084__vss n1086__vss 48.49e-3
rk4839 n1086__vss n1087__vss 187.7e-3
rk4840 n1087__vss n1088__vss 290.3e-3
rk4841 n1087__vss n1089__vss 103e-3
rk4842 n1089__vss n1090__vss 75.4253
rk4843 n1088__vss n1051__vss 322.9e-3
rk4844 n1089__vss n1091__vss 571.3e-3
rk4845 n1091__vss n1092__vss 75.4386
rk4846 n1091__vss n1093__vss 628.3e-3
rk4847 n1093__vss n1094__vss 19.1362
rk4848 n1093__vss n1095__vss 48.49e-3
rk4849 n1095__vss n1096__vss 242.2e-3
rk4850 n1096__vss n1097__vss 195.7e-3
rk4851 n1096__vss n1098__vss 123e-3
rk4852 n1098__vss n1099__vss 75.4138
rk4853 n1097__vss n1048__vss 227.8e-3
rk4854 n1098__vss n1100__vss 27.9e-3
rk4855 n1100__vss n1101__vss 340.1e-3
rk4856 n1101__vss n1102__vss 413.4e-3
rk4857 n1102__vss n1103__vss 191.9e-3
rk4858 n1102__vss n1104__vss 205.1e-3
rk4859 n1104__vss n1105__vss 75.408
rk4860 n1103__vss n1045__vss 223.9e-3
rk4861 n1104__vss n1106__vss 49.83e-3
rk4862 n1106__vss n1107__vss 340.1e-3
rk4863 n1107__vss n1108__vss 464.7e-3
rk4864 n1108__vss n1109__vss 185.5e-3
rk4865 n1108__vss n1110__vss 111.4e-3
rk4866 n1110__vss n1111__vss 75.4259
rk4867 n1109__vss n1042__vss 217.5e-3
rk4868 n1110__vss n1112__vss 56.62e-3
rk4869 n1112__vss n1113__vss 357.6e-3
rk4870 n1113__vss n1114__vss 75.1686
rk4871 n1113__vss n1115__vss 102e-3
rk4872 n1115__vss n1116__vss 558.4e-3
rk4873 n1116__vss n1117__vss 411.3e-3
rk4874 n1117__vss n1118__vss 185.5e-3
rk4875 n1117__vss n1119__vss 157.5e-3
rk4876 n1119__vss n1120__vss 75.4259
rk4877 n1118__vss n1038__vss 217.5e-3
rk4878 n1119__vss n1121__vss 56.62e-3
rk4879 n1121__vss n1122__vss 357.6e-3
rk4880 n1122__vss n1123__vss 75.1686
rk4881 n1122__vss n1124__vss 102e-3
rk4882 n1124__vss n1125__vss 558.4e-3
rk4883 n1125__vss n1126__vss 388.6e-3
rk4884 n1126__vss n1127__vss 192.5e-3
rk4885 n1126__vss n1128__vss 197.6e-3
rk4886 n1128__vss n1129__vss 75.3578
rk4887 n1127__vss n1034__vss 226.5e-3
rk4888 n1128__vss n1130__vss 175.4e-3
rk4889 n1130__vss n1131__vss 29.59e-3
rk4890 n1131__vss n1132__vss 75.3611
rk4891 n1131__vss n1133__vss 347.7e-3
rk4892 n1133__vss n1134__vss 75.418
rk4893 n1133__vss n1135__vss 324.8e-3
rk4894 n1135__vss n1136__vss 520.2e-3
rk4895 n1136__vss n1137__vss 183.5e-3
rk4896 n1136__vss n1138__vss 140.9e-3
rk4897 n1138__vss n1139__vss 37.8441
rk4898 n1137__vss n1031__vss 213.4e-3
rk4899 n1138__vss n1140__vss 467.3e-3
rk4900 n1140__vss n1141__vss 132.1e-3
rk4901 n1141__vss n1142__vss 37.8504
rk4902 n1141__vss n1143__vss 619.1e-3
rk4903 n1143__vss n1144__vss 19.1741
rk4904 n1143__vss n1145__vss 303.5e-3
rk4905 n1145__vss n1146__vss 75.418
rk4906 n1145__vss n1147__vss 240.4e-3
rk4907 n1147__vss n1148__vss 184e-3
rk4908 n1147__vss n1149__vss 85.77e-3
rk4909 n1149__vss n1150__vss 578.4e-3
rk4910 n1150__vss n1151__vss 184e-3
rk4911 n1148__vss n1028__vss 214.9e-3
rk4912 n1150__vss n1152__vss 82.84e-3
rk4913 n1152__vss n1153__vss 37.8441
rk4914 n1151__vss n1025__vss 214.9e-3
rk4915 n1152__vss n1154__vss 467.3e-3
rk4916 n1154__vss n1155__vss 132.1e-3
rk4917 n1155__vss n1156__vss 37.8504
rk4918 n1155__vss n1157__vss 619.1e-3
rk4919 n1157__vss n1158__vss 19.1741
rk4920 n1157__vss n1159__vss 198e-3
rk4921 n1159__vss n1160__vss 184.2e-3
rk4922 n1159__vss n1161__vss 84.09e-3
rk4923 n1161__vss n1162__vss 75.4595
rk4924 n1160__vss n1022__vss 216.3e-3
rk4925 n1161__vss n1163__vss 353.4e-3
rk4926 n1163__vss n1164__vss 660e-3
rk4927 n1164__vss n1165__vss 37.8441
rk4928 n1164__vss n1166__vss 467.3e-3
rk4929 n1166__vss n1167__vss 75.76e-3
rk4930 n1167__vss n1168__vss 184e-3
rk4931 n1167__vss n1169__vss 57.83e-3
rk4932 n1169__vss n1170__vss 37.8504
rk4933 n1168__vss n1019__vss 214.9e-3
rk4934 n1169__vss n1171__vss 619.1e-3
rk4935 n1171__vss n1172__vss 19.1741
rk4936 n1171__vss n1173__vss 214.1e-3
rk4937 n1173__vss n1174__vss 242.6e-3
rk4938 n1173__vss n1175__vss 62.12e-3
rk4939 n1175__vss n1176__vss 37.8279
rk4940 n1174__vss n1017__vss 167.3e-3
rk4941 n1175__vss n1177__vss 245.4e-3
rk4942 n1177__vss n1178__vss 48.49e-3
rk4943 n1178__vss n1179__vss 37.8274
rk4944 n1178__vss n1180__vss 209.8e-3
rk4945 n1180__vss n1181__vss 37.827
rk4946 n1180__vss n1182__vss 395.4e-3
rk4947 n1182__vss n1183__vss 90.02e-3
rk4948 n1183__vss n1184__vss 75.2497
rk4949 n1182__vss n1185__vss 2.7809
rk4950 n1185__vss n1186__vss 158.7e-3
rk4951 n1186__vss n1187__vss 58.74e-3
rk4952 n1187__vss n1188__vss 209.8e-3
rk4953 n1188__vss n1189__vss 416.5e-3
rk4954 n1189__vss n1190__vss 30.55e-3
rk4955 n1190__vss n1191__vss 179.2e-3
rk4956 n1191__vss n1192__vss 442.7e-3
rk4957 n1183__vss n1193__vss 75.1478
rk4958 n1183__vss n1194__vss 75.2536
rk4959 n1185__vss n1195__vss 37.8519
rk4960 n1187__vss n1196__vss 75.3645
rk4961 n1188__vss n1197__vss 75.3645
rk4962 n1189__vss n1198__vss 75.3637
rk4963 n1191__vss n1199__vss 75.3578
rk4964 n1192__vss n1200__vss 639.4e-3
rk4965 n1200__vss n1201__vss 135.6e-3
rk4966 n1201__vss n1202__vss 479.1e-3
rk4967 n1202__vss n1203__vss 488.9e-3
rk4968 n1203__vss n1204__vss 30.55e-3
rk4969 n1204__vss n1205__vss 179.2e-3
rk4970 n1205__vss n1206__vss 442.7e-3
rk4971 n1192__vss n1207__vss 19.1261
rk4972 n1200__vss n1208__vss 37.853
rk4973 n1202__vss n1209__vss 37.8467
rk4974 n1203__vss n1210__vss 75.3637
rk4975 n1205__vss n1211__vss 75.368
rk4976 n1206__vss n1212__vss 639.4e-3
rk4977 n1212__vss n1213__vss 135.6e-3
rk4978 n1213__vss n1214__vss 479.1e-3
rk4979 n1214__vss n1215__vss 455.4e-3
rk4980 n1215__vss n1216__vss 30.55e-3
rk4981 n1216__vss n1217__vss 179.2e-3
rk4982 n1217__vss n702__vss 279.7e-3
rk4983 n1206__vss n1218__vss 19.1261
rk4984 n1212__vss n1219__vss 37.853
rk4985 n1214__vss n1220__vss 37.8467
rk4986 n1215__vss n1221__vss 75.3637
rk4987 n1217__vss n1222__vss 75.3578
rk4988 n702__vss n645__vss 236.9e-3
rk4989 n645__vss n1223__vss 151.1e-3
rk4990 n1223__vss n633__vss 32e-3
rk4991 n633__vss n1224__vss 164.4e-3
rk4992 n1224__vss n1225__vss 209.8e-3
rk4993 n1225__vss n1226__vss 322e-3
rk4994 n1226__vss n1227__vss 50.83e-3
rk4995 n1227__vss n1228__vss 412.3e-3
rk4996 n1228__vss n1229__vss 351.9e-3
rk4997 n1229__vss n1230__vss 338.5e-3
rk4998 n1230__vss n1231__vss 506.8e-3
rk4999 n1231__vss n1232__vss 54.24e-3
rk5000 n1232__vss n1233__vss 527.5e-3
rk5001 n1233__vss n1234__vss 340.1e-3
rk5002 n1234__vss n1235__vss 44.21e-3
rk5003 n1235__vss n1236__vss 533.3e-3
rk5004 n1236__vss n1237__vss 340.1e-3
rk5005 n1237__vss n1238__vss 48.92e-3
rk5006 n1238__vss n1239__vss 628.4e-3
rk5007 n1239__vss n1240__vss 558.4e-3
rk5008 n1240__vss n1241__vss 102e-3
rk5009 n1241__vss n1242__vss 357.6e-3
rk5010 n1242__vss n1243__vss 49.63e-3
rk5011 n1243__vss n1244__vss 589.6e-3
rk5012 n1244__vss n1245__vss 340.1e-3
rk5013 n1245__vss n1246__vss 55.78e-3
rk5014 n1246__vss n1247__vss 640.9e-3
rk5015 n1247__vss n1248__vss 340.1e-3
rk5016 n1248__vss n1249__vss 49.83e-3
rk5017 n1249__vss n1250__vss 338.7e-3
rk5018 n1250__vss n1251__vss 47.1e-3
rk5019 n1251__vss n1252__vss 625.1e-3
rk5020 n1252__vss n1253__vss 571.3e-3
rk5021 n1253__vss n1254__vss 289.4e-3
rk5022 n1254__vss n1255__vss 48.49e-3
rk5023 n1255__vss n1256__vss 628.3e-3
rk5024 n1256__vss n1257__vss 571.3e-3
rk5025 n1257__vss n1258__vss 274e-3
rk5026 n1258__vss n1259__vss 48.49e-3
rk5027 n1259__vss n1260__vss 628.3e-3
rk5028 n1260__vss n1261__vss 571.3e-3
rk5029 n1261__vss n1262__vss 289.4e-3
rk5030 n1262__vss n1263__vss 48.49e-3
rk5031 n1263__vss n1264__vss 628.3e-3
rk5032 n1264__vss n1265__vss 672.8e-3
rk5033 n1265__vss n1266__vss 147.4e-3
rk5034 n1266__vss n1267__vss 75.4606
rk5035 n1224__vss n1268__vss 37.827
rk5036 n1225__vss n1269__vss 37.8273
rk5037 n1227__vss n1270__vss 75.3993
rk5038 n1228__vss n1271__vss 75.1418
rk5039 n1230__vss n1272__vss 75.1418
rk5040 n1232__vss n1273__vss 75.4022
rk5041 n1235__vss n1274__vss 75.4528
rk5042 n1238__vss n1275__vss 75.4487
rk5043 n1241__vss n1276__vss 75.1686
rk5044 n1243__vss n1277__vss 75.4533
rk5045 n1246__vss n1278__vss 75.4539
rk5046 n1249__vss n1279__vss 75.408
rk5047 n1251__vss n1280__vss 19.1336
rk5048 n1252__vss n1281__vss 75.4386
rk5049 n1253__vss n1282__vss 75.4253
rk5050 n1255__vss n1283__vss 19.1362
rk5051 n1256__vss n1284__vss 75.4386
rk5052 n1257__vss n1285__vss 75.4253
rk5053 n1259__vss n1286__vss 19.1362
rk5054 n1260__vss n1287__vss 75.4386
rk5055 n1261__vss n1288__vss 75.4253
rk5056 n1263__vss n1289__vss 19.1362
rk5057 n1264__vss n1290__vss 75.4386
rk5058 n1265__vss n1291__vss 75.4748
rk5059 n1013__vss n1014__vss 4.1333
rk5060 n913__vss n1015__vss 16.67e-3
rk5061 n1013__vss n1016__vss 1.0333
rk5062 n919__vss n1017__vss 8.333e-3
rk5063 n1013__vss n1018__vss 1.0333
rk5064 n926__vss n1020__vss 8.333e-3
rk5065 n1013__vss n1021__vss 1.0333
rk5066 n934__vss n1023__vss 8.333e-3
rk5067 n1013__vss n1024__vss 1.0333
rk5068 n939__vss n1026__vss 8.333e-3
rk5069 n1013__vss n1027__vss 1.0333
rk5070 n1013__vss n1029__vss 1.0333
rk5071 n944__vss n1030__vss 8.333e-3
rk5072 n1013__vss n1031__vss 1.0333
rk5073 n949__vss n1032__vss 8.333e-3
rk5074 n1013__vss n1033__vss 1.0333
rk5075 n954__vss n1035__vss 8.333e-3
rk5076 n1013__vss n1036__vss 1.0333
rk5077 n960__vss n1037__vss 8.333e-3
rk5078 n1013__vss n1039__vss 1.0333
rk5079 n966__vss n1040__vss 8.333e-3
rk5080 n1013__vss n1041__vss 1.0333
rk5081 n971__vss n1043__vss 8.333e-3
rk5082 n1013__vss n1044__vss 1.0333
rk5083 n1013__vss n1046__vss 1.0333
rk5084 n978__vss n1047__vss 8.333e-3
rk5085 n1013__vss n1049__vss 1.0333
rk5086 n986__vss n1050__vss 8.333e-3
rk5087 n1013__vss n1052__vss 1.0333
rk5088 n991__vss n1053__vss 8.333e-3
rk5089 n1013__vss n1054__vss 1.0333
rk5090 n997__vss n1055__vss 8.333e-3
rk5091 n1013__vss n1056__vss 1.0333
rk5092 n1004__vss n1058__vss 8.333e-3
rk5093 n1013__vss n1059__vss 1.0333
rk5094 n1010__vss n1060__vss 8.333e-3
rk5095 n1013__vss n1062__vss 31
rk5096 n1013__vss n1064__vss 3.1
rk5097 n1013__vss n1066__vss 20.6667
rk5098 n1013__vss n1073__vss 3.1
rk5099 n1013__vss n1077__vss 31
rk5100 n1013__vss n1082__vss 3.1
rk5101 n1013__vss n1086__vss 31
rk5102 n1013__vss n1091__vss 3.1
rk5103 n1013__vss n1095__vss 31
rk5104 n1013__vss n1100__vss 20.6667
rk5105 n1013__vss n1101__vss 6.2
rk5106 n1013__vss n1106__vss 20.6667
rk5107 n1013__vss n1107__vss 6.2
rk5108 n1013__vss n1112__vss 20.6667
rk5109 n1013__vss n1115__vss 6.2
rk5110 n1013__vss n1116__vss 6.2
rk5111 n1013__vss n1121__vss 20.6667
rk5112 n1013__vss n1124__vss 6.2
rk5113 n1013__vss n1125__vss 6.2
rk5114 n1013__vss n1130__vss 7.75
rk5115 n1013__vss n1135__vss 5.1667
rk5116 n1013__vss n1140__vss 3.1
rk5117 n1013__vss n1143__vss 12.4
rk5118 n1013__vss n1149__vss 5.1667
rk5119 n1013__vss n1154__vss 3.1
rk5120 n1013__vss n1157__vss 12.4
rk5121 n1013__vss n1163__vss 5.1667
rk5122 n1013__vss n1166__vss 3.1
rk5123 n1013__vss n1171__vss 12.4
rk5124 n1013__vss n1177__vss 6.2
rk5125 n1013__vss n1182__vss 7.75
rk5126 n1013__vss n1186__vss 6.2
rk5127 n1013__vss n1190__vss 7.75
rk5128 n1013__vss n1192__vss 12.4
rk5129 n1013__vss n1201__vss 3.1
rk5130 n1013__vss n1204__vss 7.75
rk5131 n1013__vss n1206__vss 12.4
rk5132 n1013__vss n1213__vss 3.1
rk5133 n1013__vss n1216__vss 7.75
rk5134 n1013__vss n1223__vss 4.1333
rk5135 n1013__vss n1226__vss 20.6667
rk5136 n1013__vss n1229__vss 4.4286
rk5137 n1013__vss n1231__vss 20.6667
rk5138 n1013__vss n1233__vss 6.2
rk5139 n1013__vss n1234__vss 20.6667
rk5140 n1013__vss n1236__vss 6.2
rk5141 n1013__vss n1237__vss 20.6667
rk5142 n1013__vss n1239__vss 6.2
rk5143 n1013__vss n1240__vss 6.2
rk5144 n1013__vss n1242__vss 20.6667
rk5145 n1013__vss n1244__vss 6.2
rk5146 n1013__vss n1245__vss 20.6667
rk5147 n1013__vss n1247__vss 6.2
rk5148 n1013__vss n1248__vss 20.6667
rk5149 n1013__vss n1250__vss 31
rk5150 n1013__vss n1252__vss 3.1
rk5151 n1013__vss n1254__vss 31
rk5152 n1013__vss n1256__vss 3.1
rk5153 n1013__vss n1258__vss 31
rk5154 n1013__vss n1260__vss 3.1
rk5155 n1013__vss n1262__vss 31
rk5156 n1013__vss n1264__vss 3.1
rk5157 n1013__vss n1266__vss 20.6667
rk5158 n230__i1__net2 n231__i1__net2 323.1e-3
rk5159 n231__i1__net2 n233__i1__net2 148.3e-3
rk5160 n230__i1__net2 n232__i1__net2 5.2293
rk5161 n233__i1__net2 n234__i1__net2 271.8e-3
rk5162 n232__i1__net2 n233__i1__net2 3.1
rk5163 n235__i1__net2 n236__i1__net2 75.293
rk5164 n236__i1__net2 n237__i1__net2 69.31e-3
rk5165 n237__i1__net2 n238__i1__net2 351.9e-3
rk5166 n235__i1__net2 n237__i1__net2 3.75
rk5167 i1__net3 n2__i1__net3 15.125
rk5169 n5__i1__net3 n6__i1__net3 8.857e-3
rk5171 n4__i1__net3 n5__i1__net3 7.75
rk5172 n4__i1__i13__net1 n61__i1__i13__net1 125e-3
rk5173 n2__i1__i13__net1 n62__i1__i13__net1 125e-3
rk5174 n2__i1__i12__net1 n29__i1__i12__net1 125e-3
rk5175 n4__i1__i12__net1 n30__i1__i12__net1 125e-3
rk5176 n1678__vddio n1680__vddio 187.3e-3
rk5177 n1680__vddio n1681__vddio 231e-3
rk5178 n1681__vddio n1682__vddio 316.2e-3
rk5179 n1682__vddio n1683__vddio 27.62e-3
rk5180 n1683__vddio n1684__vddio 332.4e-3
rk5181 n1679__vddio n1680__vddio 5.1667
rk5182 n1679__vddio n1682__vddio 3.1
rk5183 n1292__vss n1294__vss 44.28e-3
rk5184 n1294__vss n1295__vss 121.7e-3
rk5185 n1295__vss n1296__vss 240.5e-3
rk5186 n1296__vss n1297__vss 103.3e-3
rk5188 n1293__vss n1294__vss 75
rk5189 n1293__vss n1296__vss 3.75
rk5192 n6__i1__i12__net1 n33__i1__i12__net1 125e-3
rk5193 n8__i1__i12__net1 n34__i1__i12__net1 125e-3
rk5194 n239__i1__net2 n240__i1__net2 75.293
rk5195 n240__i1__net2 n241__i1__net2 69.31e-3
rk5196 n241__i1__net2 n242__i1__net2 351.9e-3
rk5197 n239__i1__net2 n241__i1__net2 3.75
rk5198 n243__i1__net2 n244__i1__net2 323.1e-3
rk5199 n244__i1__net2 n246__i1__net2 148.3e-3
rk5200 n243__i1__net2 n245__i1__net2 5.2293
rk5201 n246__i1__net2 n247__i1__net2 271.8e-3
rk5202 n245__i1__net2 n246__i1__net2 3.1
rk5203 n8__i1__net3 n10__i1__net3 25.45e-3
rk5204 n9__i1__net3 n10__i1__net3 15
rk5206 n13__i1__net3 n14__i1__net3 8.139e-3
rk5208 n12__i1__net3 n13__i1__net3 7.75
rk5209 n12__i1__i13__net1 n73__i1__i13__net1 125e-3
rk5210 n10__i1__i13__net1 n74__i1__i13__net1 125e-3
rk5211 n10__i1__i12__net1 n37__i1__i12__net1 125e-3
rk5212 n12__i1__i12__net1 n38__i1__i12__net1 125e-3
rk5213 n1299__vss n1301__vss 240.5e-3
rk5214 n1299__vss n1302__vss 115.4e-3
rk5215 n1302__vss n1303__vss 171.4e-3
rk5216 n1301__vss n1304__vss 185.5e-3
rk5217 n1300__vss n1301__vss 3.75
rk5218 n1300__vss n1302__vss 75
rk5219 n1685__vddio n1687__vddio 187.3e-3
rk5220 n1687__vddio n1688__vddio 231e-3
rk5221 n1688__vddio n1689__vddio 316.2e-3
rk5222 n1689__vddio n1690__vddio 27.62e-3
rk5223 n1690__vddio n1691__vddio 332.4e-3
rk5224 n1686__vddio n1687__vddio 5.1667
rk5225 n1686__vddio n1689__vddio 3.1
rk5226 n16__i1__i13__net1 n85__i1__i13__net1 125e-3
rk5227 n14__i1__i13__net1 n86__i1__i13__net1 125e-3
rk5228 n14__i1__i12__net1 n41__i1__i12__net1 125e-3
rk5229 n16__i1__i12__net1 n42__i1__i12__net1 125e-3
rk5230 n248__i1__net2 n249__i1__net2 323.1e-3
rk5231 n249__i1__net2 n251__i1__net2 148.3e-3
rk5232 n248__i1__net2 n250__i1__net2 5.2293
rk5233 n251__i1__net2 n252__i1__net2 271.8e-3
rk5234 n250__i1__net2 n251__i1__net2 3.1
rk5235 n253__i1__net2 n254__i1__net2 75.293
rk5236 n254__i1__net2 n255__i1__net2 69.31e-3
rk5237 n255__i1__net2 n256__i1__net2 351.9e-3
rk5238 n253__i1__net2 n255__i1__net2 3.75
rk5239 n16__i1__net3 n17__i1__net3 15.126
rk5241 n20__i1__net3 n21__i1__net3 5.905e-3
rk5243 n19__i1__net3 n20__i1__net3 7.75
rk5246 n18__i1__i12__net1 n45__i1__i12__net1 125e-3
rk5247 n20__i1__i12__net1 n46__i1__i12__net1 125e-3
rk5248 n1692__vddio n1694__vddio 187.3e-3
rk5249 n1694__vddio n1695__vddio 231e-3
rk5250 n1695__vddio n1696__vddio 316.2e-3
rk5251 n1696__vddio n1697__vddio 27.62e-3
rk5252 n1697__vddio n1698__vddio 330.7e-3
rk5253 n1693__vddio n1694__vddio 5.1667
rk5254 n1693__vddio n1696__vddio 3.1
rk5255 n1306__vss n1308__vss 240.5e-3
rk5256 n1306__vss n1309__vss 117.9e-3
rk5257 n1309__vss n1310__vss 168.7e-3
rk5258 n1308__vss n1311__vss 185.5e-3
rk5259 n1307__vss n1308__vss 3.75
rk5260 n1307__vss n1309__vss 75
rk5261 n24__i1__i13__net1 n101__i1__i13__net1 125e-3
rk5262 n22__i1__i13__net1 n102__i1__i13__net1 125e-3
rk5263 n22__i1__i12__net1 n49__i1__i12__net1 125e-3
rk5264 n24__i1__i12__net1 n50__i1__i12__net1 125e-3
rk5265 n257__i1__net2 n258__i1__net2 323.1e-3
rk5266 n258__i1__net2 n260__i1__net2 148.3e-3
rk5267 n257__i1__net2 n259__i1__net2 5.2293
rk5268 n260__i1__net2 n261__i1__net2 271.8e-3
rk5269 n259__i1__net2 n260__i1__net2 3.1
rk5270 n262__i1__net2 n263__i1__net2 75.293
rk5271 n263__i1__net2 n264__i1__net2 69.31e-3
rk5272 n264__i1__net2 n265__i1__net2 351.9e-3
rk5273 n262__i1__net2 n264__i1__net2 3.75
rk5275 n25__i1__net3 n26__i1__net3 8.857e-3
rk5277 n24__i1__net3 n25__i1__net3 7.75
rk5278 n28__i1__net3 n29__i1__net3 15.125
rk5283 n1699__vddio n1701__vddio 187.3e-3
rk5284 n1701__vddio n1702__vddio 231e-3
rk5285 n1702__vddio n1703__vddio 316.2e-3
rk5286 n1703__vddio n1704__vddio 27.62e-3
rk5287 n1704__vddio n1705__vddio 332.4e-3
rk5288 n1700__vddio n1701__vddio 5.1667
rk5289 n1700__vddio n1703__vddio 3.1
rk5290 n1554__vss n1555__vss 121.7e-3
rk5291 n1555__vss n1556__vss 240.5e-3
rk5292 n1556__vss n1557__vss 103.3e-3
rk5294 n1554__vss n1559__vss 172.2e-3
rk5295 n1553__vss n1554__vss 75
rk5296 n1553__vss n1556__vss 3.75
rk5299 n266__i1__net2 n267__i1__net2 323.1e-3
rk5300 n267__i1__net2 n269__i1__net2 148.3e-3
rk5301 n266__i1__net2 n268__i1__net2 5.2293
rk5302 n269__i1__net2 n270__i1__net2 271.8e-3
rk5303 n268__i1__net2 n269__i1__net2 3.1
rk5304 n271__i1__net2 n272__i1__net2 75.293
rk5305 n272__i1__net2 n273__i1__net2 69.31e-3
rk5306 n273__i1__net2 n274__i1__net2 351.9e-3
rk5307 n271__i1__net2 n273__i1__net2 3.75
rk5308 n35__i1__i13__net1 n113__i1__i13__net1 125e-3
rk5309 n34__i1__i13__net1 n114__i1__i13__net1 125e-3
rk5310 n1706__vddio n1707__vddio 459.3e-3
rk5311 n1707__vddio n1709__vddio 27.62e-3
rk5312 n1709__vddio n1710__vddio 316.2e-3
rk5313 n1710__vddio n1711__vddio 231e-3
rk5314 n1711__vddio n1712__vddio 187.3e-3
rk5315 n1708__vddio n1709__vddio 3.1
rk5316 n1708__vddio n1711__vddio 5.1667
rk5317 n1560__vss n1562__vss 117.9e-3
rk5318 n1562__vss n1563__vss 84.83e-3
rk5319 n1560__vss n1564__vss 240.5e-3
rk5320 n1564__vss n1565__vss 185.5e-3
rk5321 n1561__vss n1562__vss 75
rk5322 n1561__vss n1564__vss 3.75
rk5323 n40__i1__i13__net1 n117__i1__i13__net1 125e-3
rk5324 n38__i1__i13__net1 n118__i1__i13__net1 125e-3
rk5325 n2__i1__net4 n13__i1__net4 125e-3
rk5326 n4__i1__net4 n14__i1__net4 125e-3
rk5327 n275__i1__net2 n276__i1__net2 323.1e-3
rk5328 n276__i1__net2 n278__i1__net2 148.3e-3
rk5329 n275__i1__net2 n277__i1__net2 5.2293
rk5330 n278__i1__net2 n279__i1__net2 271.8e-3
rk5331 n277__i1__net2 n278__i1__net2 3.1
rk5332 n280__i1__net2 n281__i1__net2 75.293
rk5333 n281__i1__net2 n282__i1__net2 69.31e-3
rk5334 n282__i1__net2 n283__i1__net2 351.9e-3
rk5335 n280__i1__net2 n282__i1__net2 3.75
rk5337 n63__i1__i12__net1 n64__i1__i12__net1 148.6e-3
rk5338 n62__i1__i12__net1 n63__i1__i12__net1 7.75
rk5339 n65__i1__i12__net1 n66__i1__i12__net1 15.125
rk5340 n43__i1__i13__net1 n125__i1__i13__net1 125e-3
rk5341 n42__i1__i13__net1 n126__i1__i13__net1 125e-3
rk5342 n1713__vddio n1715__vddio 187.3e-3
rk5343 n1715__vddio n1716__vddio 231e-3
rk5344 n1716__vddio n1717__vddio 316.2e-3
rk5345 n1717__vddio n1718__vddio 27.62e-3
rk5346 n1718__vddio n1719__vddio 327.7e-3
rk5347 n1714__vddio n1715__vddio 5.1667
rk5348 n1714__vddio n1717__vddio 3.1
rk5349 n1566__vss n1568__vss 240.5e-3
rk5350 n1566__vss n1569__vss 117.9e-3
rk5351 n1569__vss n1570__vss 171.7e-3
rk5352 n1568__vss n1571__vss 185.5e-3
rk5353 n1567__vss n1568__vss 3.75
rk5354 n1567__vss n1569__vss 75
rk5355 n6__i1__net4 n17__i1__net4 125e-3
rk5356 n8__i1__net4 n18__i1__net4 125e-3
rk5357 n48__i1__i13__net1 n129__i1__i13__net1 125e-3
rk5358 n46__i1__i13__net1 n130__i1__i13__net1 125e-3
rk5359 n1572__vss n1573__vss 15.2439
rk5360 n1573__vss n1574__vss 21.14e-3
rk5361 n1574__vss n1575__vss 87.08e-3
rk5362 n1575__vss n1576__vss 78.17e-3
rk5363 n1576__vss n1577__vss 49.94e-3
rk5364 n1577__vss n1578__vss 21.14e-3
rk5365 n1578__vss n1579__vss 15.2735
rk5366 n1574__vss n1580__vss 15.2142
rk5367 n1575__vss n1581__vss 15.1676
rk5368 n1576__vss n1582__vss 15.1708
rk5369 n1578__vss n1583__vss 15.2204
rk5370 n1013__vss n1574__vss 2.0667
rk5371 n1013__vss n1578__vss 1.55
rk5372 n284__i1__net2 n285__i1__net2 323.1e-3
rk5373 n285__i1__net2 n287__i1__net2 148.3e-3
rk5374 n284__i1__net2 n286__i1__net2 5.2293
rk5375 n287__i1__net2 n288__i1__net2 271.8e-3
rk5376 n286__i1__net2 n287__i1__net2 3.1
rk5377 n289__i1__net2 n290__i1__net2 75.293
rk5378 n290__i1__net2 n291__i1__net2 69.31e-3
rk5379 n291__i1__net2 n292__i1__net2 351.9e-3
rk5380 n289__i1__net2 n291__i1__net2 3.75
rk5381 n51__i1__i13__net1 n133__i1__i13__net1 125e-3
rk5382 n50__i1__i13__net1 n134__i1__i13__net1 125e-3
rk5383 n1738__vddio n1740__vddio 187.3e-3
rk5384 n1740__vddio n1741__vddio 231e-3
rk5385 n1741__vddio n1742__vddio 316.2e-3
rk5386 n1742__vddio n1743__vddio 27.62e-3
rk5387 n1743__vddio n1744__vddio 332.4e-3
rk5388 n1739__vddio n1740__vddio 5.1667
rk5389 n1739__vddio n1742__vddio 3.1
rk5390 n1587__vss n1589__vss 44.28e-3
rk5391 n1589__vss n1590__vss 121.7e-3
rk5392 n1590__vss n1591__vss 240.5e-3
rk5393 n1591__vss n1592__vss 103.3e-3
rk5395 n1588__vss n1589__vss 75
rk5396 n1588__vss n1591__vss 3.75
rk5397 n56__i1__i13__net1 n137__i1__i13__net1 125e-3
rk5398 n54__i1__i13__net1 n138__i1__i13__net1 125e-3
rk5399 n23__piso_out n28__piso_out 250e-3
rk5400 n9__i1__net4 n22__i1__net4 250e-3
rk5401 n293__i1__net2 n294__i1__net2 323.1e-3
rk5402 n294__i1__net2 n296__i1__net2 148.3e-3
rk5403 n293__i1__net2 n295__i1__net2 5.2293
rk5404 n296__i1__net2 n297__i1__net2 271.8e-3
rk5405 n295__i1__net2 n296__i1__net2 3.1
rk5406 n298__i1__net2 n299__i1__net2 75.293
rk5407 n299__i1__net2 n300__i1__net2 69.31e-3
rk5408 n300__i1__net2 n301__i1__net2 351.9e-3
rk5409 n298__i1__net2 n300__i1__net2 3.75
rk5410 n59__i1__i13__net1 n141__i1__i13__net1 125e-3
rk5411 n58__i1__i13__net1 n142__i1__i13__net1 125e-3
rk5412 n24__piso_out n31__piso_out 250e-3
rk5413 n1745__vddio n1747__vddio 187.3e-3
rk5414 n1747__vddio n1748__vddio 231e-3
rk5415 n1748__vddio n1749__vddio 316.2e-3
rk5416 n1749__vddio n1750__vddio 27.62e-3
rk5417 n1750__vddio n1751__vddio 327.7e-3
rk5418 n1746__vddio n1747__vddio 5.1667
rk5419 n1746__vddio n1749__vddio 3.1
rk5420 n1595__vss n1596__vss 121.7e-3
rk5421 n1596__vss n1597__vss 240.5e-3
rk5422 n1597__vss n1598__vss 103.3e-3
rk5424 n1595__vss n1600__vss 172.2e-3
rk5425 n1594__vss n1595__vss 75
rk5426 n1594__vss n1597__vss 3.75
rk5427 n11__i1__net4 n23__i1__net4 250e-3
rk5428 n5__i1__i11__outinv n6__i1__i11__outinv 15.2961
rk5429 n6__i1__i11__outinv n7__i1__i11__outinv 132.2e-3
rk5430 n6__i1__i11__outinv n8__i1__i11__outinv 31.2241
rk5431 n7__i1__i11__outinv n9__i1__i11__outinv 15.2128
rk5435 n302__i1__net2 n303__i1__net2 323.1e-3
rk5436 n303__i1__net2 n305__i1__net2 148.3e-3
rk5437 n302__i1__net2 n304__i1__net2 5.2293
rk5438 n305__i1__net2 n306__i1__net2 271.8e-3
rk5439 n304__i1__net2 n305__i1__net2 3.1
rk5440 n307__i1__net2 n308__i1__net2 75.293
rk5441 n308__i1__net2 n309__i1__net2 69.31e-3
rk5442 n309__i1__net2 n310__i1__net2 351.9e-3
rk5443 n307__i1__net2 n309__i1__net2 3.75
rk5444 n79__i1__i13__net1 n149__i1__i13__net1 125e-3
rk5445 n78__i1__i13__net1 n150__i1__i13__net1 125e-3
rk5446 n1752__vddio n1754__vddio 187.3e-3
rk5447 n1754__vddio n1755__vddio 231e-3
rk5448 n1755__vddio n1756__vddio 316.2e-3
rk5449 n1756__vddio n1757__vddio 27.62e-3
rk5450 n1757__vddio n1758__vddio 332.4e-3
rk5451 n1753__vddio n1754__vddio 5.1667
rk5452 n1753__vddio n1756__vddio 3.1
rk5453 n1601__vss n1603__vss 117.9e-3
rk5454 n1603__vss n1604__vss 84.83e-3
rk5455 n1601__vss n1605__vss 240.5e-3
rk5456 n1605__vss n1606__vss 185.5e-3
rk5457 n1602__vss n1603__vss 75
rk5458 n1602__vss n1605__vss 3.75
rk5459 n84__i1__i13__net1 n151__i1__i13__net1 125e-3
rk5460 n82__i1__i13__net1 n152__i1__i13__net1 125e-3
rk5461 n311__i1__net2 n312__i1__net2 75.293
rk5462 n312__i1__net2 n313__i1__net2 69.31e-3
rk5463 n313__i1__net2 n314__i1__net2 351.9e-3
rk5464 n311__i1__net2 n313__i1__net2 3.75
rk5465 n9__piso_outinv n15__piso_outinv 250e-3
rk5466 n315__i1__net2 n316__i1__net2 323.1e-3
rk5467 n316__i1__net2 n318__i1__net2 148.3e-3
rk5468 n315__i1__net2 n317__i1__net2 5.2293
rk5469 n318__i1__net2 n319__i1__net2 271.8e-3
rk5470 n317__i1__net2 n318__i1__net2 3.1
rk5471 n91__i1__i13__net1 n153__i1__i13__net1 125e-3
rk5472 n90__i1__i13__net1 n154__i1__i13__net1 125e-3
rk5473 i1__i11__outinv n10__i1__i11__outinv 250e-3
rk5474 n1607__vss n1609__vss 185.5e-3
rk5475 n1609__vss n1610__vss 240.5e-3
rk5476 n1610__vss n1611__vss 117.9e-3
rk5477 n1611__vss n1612__vss 171.7e-3
rk5478 n1608__vss n1609__vss 3.75
rk5479 n1608__vss n1611__vss 75
rk5480 n1759__vddio n1761__vddio 187.3e-3
rk5481 n1761__vddio n1762__vddio 231e-3
rk5482 n1762__vddio n1763__vddio 316.2e-3
rk5483 n1763__vddio n1764__vddio 27.62e-3
rk5484 n1764__vddio n1765__vddio 326.2e-3
rk5485 n1760__vddio n1761__vddio 5.1667
rk5486 n1760__vddio n1763__vddio 3.1
rk5487 n11__piso_outinv n16__piso_outinv 250e-3
rk5488 n100__i1__i13__net1 n155__i1__i13__net1 125e-3
rk5489 n98__i1__i13__net1 n156__i1__i13__net1 125e-3
rk5490 n24__i1__net4 n25__i1__net4 15.4801
rk5491 n25__i1__net4 n26__i1__net4 31.2379
rk5492 n25__i1__net4 n27__i1__net4 15.2315
rk5493 n320__i1__net2 n321__i1__net2 75.293
rk5494 n321__i1__net2 n322__i1__net2 69.31e-3
rk5495 n322__i1__net2 n323__i1__net2 351.9e-3
rk5496 n320__i1__net2 n322__i1__net2 3.75
rk5497 n3__i1__i11__outinv n11__i1__i11__outinv 250e-3
rk5498 n13__piso_outinv n17__piso_outinv 250e-3
rk5499 n324__i1__net2 n325__i1__net2 323.1e-3
rk5500 n325__i1__net2 n327__i1__net2 148.3e-3
rk5501 n324__i1__net2 n326__i1__net2 5.2293
rk5502 n327__i1__net2 n328__i1__net2 271.8e-3
rk5503 n326__i1__net2 n327__i1__net2 3.1
rk5504 n123__i1__i13__net1 n157__i1__i13__net1 125e-3
rk5505 n122__i1__i13__net1 n158__i1__i13__net1 125e-3
rk5506 n1766__vddio n1768__vddio 31.2196
rk5507 n1768__vddio n1769__vddio 188.8e-3
rk5508 n1769__vddio n1770__vddio 214.3e-3
rk5509 n1770__vddio n1771__vddio 413.2e-3
rk5510 n1771__vddio n1772__vddio 65.41e-3
rk5511 n1772__vddio n1773__vddio 79.86e-3
rk5512 n1773__vddio n1733__vddio 102e-3
rk5513 n1733__vddio n1774__vddio 66.03e-3
rk5514 n1774__vddio n1775__vddio 8.1268
rk5515 n1769__vddio n1776__vddio 31.1789
rk5516 n1770__vddio n1777__vddio 79.97e-3
rk5517 n1777__vddio n1778__vddio 31.3702
rk5518 n1771__vddio n1779__vddio 8.0313
rk5519 n1772__vddio n1780__vddio 8.0738
rk5520 n1773__vddio n1781__vddio 8.0371
rk5521 n1733__vddio n1782__vddio 8.0605
rk5522 n1774__vddio n1783__vddio 8.0638
rk5523 n1777__vddio n1784__vddio 31.1789
rk5524 n1767__vddio n1768__vddio 18.75
rk5525 n1767__vddio n1770__vddio 3.75
rk5526 n1730__vddio n1771__vddio 16.67e-3
rk5527 n1767__vddio n1772__vddio 2.5
rk5528 n1767__vddio n1774__vddio 1.875
rk5529 n1613__vss n1614__vss 15.3389
rk5530 n1614__vss n1615__vss 71.27e-3
rk5531 n1615__vss n1616__vss 193.5e-3
rk5532 n1616__vss n1617__vss 206.5e-3
rk5533 n1617__vss n1618__vss 61.55e-3
rk5534 n1618__vss n1619__vss 218.4e-3
rk5536 n1616__vss n1621__vss 15.263
rk5537 n1618__vss n1622__vss 15.2932
rk5538 n1619__vss n1623__vss 15.2599
rk5539 n1013__vss n1615__vss 15.5
rk5540 n1013__vss n1618__vss 3.1
rk5541 n1785__vddio n1787__vddio 187.3e-3
rk5542 n1787__vddio n1788__vddio 231e-3
rk5543 n1788__vddio n1789__vddio 316.2e-3
rk5544 n1789__vddio n1790__vddio 27.62e-3
rk5545 n1790__vddio n1791__vddio 329.1e-3
rk5546 n1786__vddio n1787__vddio 5.1667
rk5547 n1786__vddio n1789__vddio 3.1
rk5548 n1624__vss n1626__vss 44.28e-3
rk5549 n1626__vss n1627__vss 122.6e-3
rk5550 n1627__vss n1628__vss 241.4e-3
rk5551 n1628__vss n1629__vss 104.1e-3
rk5553 n1625__vss n1626__vss 75
rk5554 n1625__vss n1628__vss 3.75
rk5555 n1632__vss n1633__vss 115.8e-3
rk5556 n1633__vss n1634__vss 246.5e-3
rk5557 n1634__vss n1635__vss 97.36e-3
rk5559 n1632__vss n1637__vss 178.1e-3
rk5560 n1631__vss n1632__vss 75
rk5561 n1631__vss n1634__vss 3.75
rk5562 n1792__vddio n1793__vddio 456.3e-3
rk5563 n1793__vddio n1795__vddio 25.11e-3
rk5564 n1795__vddio n1796__vddio 318.7e-3
rk5565 n1796__vddio n1797__vddio 228e-3
rk5566 n1797__vddio n1798__vddio 190.3e-3
rk5567 n1794__vddio n1795__vddio 3.1
rk5568 n1794__vddio n1797__vddio 5.1667
rk5569 n31__i1__net3 n54__i1__net3 125e-3
rk5570 n33__i1__net3 n55__i1__net3 125e-3
rk5571 n159__i1__i13__net1 n160__i1__i13__net1 75.287
rk5572 n160__i1__i13__net1 n161__i1__i13__net1 75.22e-3
rk5573 n161__i1__i13__net1 n162__i1__i13__net1 346e-3
rk5574 n159__i1__i13__net1 n161__i1__i13__net1 3.75
rk5576 n164__i1__i13__net1 n166__i1__i13__net1 186.7e-3
rk5577 n166__i1__i13__net1 n167__i1__i13__net1 151.2e-3
rk5578 n167__i1__i13__net1 n168__i1__i13__net1 323.1e-3
rk5579 n168__i1__i13__net1 n169__i1__i13__net1 57.75e-3
rk5580 n165__i1__i13__net1 n166__i1__i13__net1 3.1
rk5581 n165__i1__i13__net1 n169__i1__i13__net1 5.1667
rk5582 n35__i1__net3 n56__i1__net3 125e-3
rk5583 n37__i1__net3 n57__i1__net3 125e-3
rk5584 n1638__vss n1640__vss 112.3e-3
rk5585 n1640__vss n1641__vss 96.14e-3
rk5586 n1638__vss n1642__vss 246.5e-3
rk5587 n1642__vss n1643__vss 179.6e-3
rk5588 n1639__vss n1640__vss 75
rk5589 n1639__vss n1642__vss 3.75
rk5590 n1799__vddio n1801__vddio 190.3e-3
rk5591 n1801__vddio n1802__vddio 228e-3
rk5592 n1802__vddio n1803__vddio 318.7e-3
rk5593 n1803__vddio n1804__vddio 25.11e-3
rk5594 n1804__vddio n1805__vddio 332.4e-3
rk5595 n1800__vddio n1801__vddio 5.1667
rk5596 n1800__vddio n1803__vddio 3.1
rk5597 n39__i1__net3 n58__i1__net3 125e-3
rk5598 n41__i1__net3 n59__i1__net3 125e-3
rk5599 n170__i1__i13__net1 n171__i1__i13__net1 75.287
rk5600 n171__i1__i13__net1 n172__i1__i13__net1 75.22e-3
rk5601 n172__i1__i13__net1 n173__i1__i13__net1 346e-3
rk5602 n170__i1__i13__net1 n172__i1__i13__net1 3.75
rk5604 n175__i1__i13__net1 n177__i1__i13__net1 186.7e-3
rk5605 n177__i1__i13__net1 n178__i1__i13__net1 151.2e-3
rk5606 n178__i1__i13__net1 n179__i1__i13__net1 323.1e-3
rk5607 n179__i1__i13__net1 n180__i1__i13__net1 57.75e-3
rk5608 n176__i1__i13__net1 n177__i1__i13__net1 3.1
rk5609 n176__i1__i13__net1 n180__i1__i13__net1 5.1667
rk5610 n43__i1__net3 n60__i1__net3 125e-3
rk5611 n45__i1__net3 n61__i1__net3 125e-3
rk5612 n1644__vss n1646__vss 115.8e-3
rk5613 n1646__vss n1647__vss 177.8e-3
rk5614 n1644__vss n1648__vss 246.5e-3
rk5615 n1648__vss n1649__vss 179.6e-3
rk5616 n1645__vss n1646__vss 75
rk5617 n1645__vss n1648__vss 3.75
rk5618 n1806__vddio n1808__vddio 190.3e-3
rk5619 n1808__vddio n1809__vddio 228e-3
rk5620 n1809__vddio n1810__vddio 318.7e-3
rk5621 n1810__vddio n1811__vddio 25.11e-3
rk5622 n1811__vddio n1812__vddio 329.5e-3
rk5623 n1807__vddio n1808__vddio 5.1667
rk5624 n1807__vddio n1810__vddio 3.1
rk5625 n47__i1__net3 n62__i1__net3 125e-3
rk5626 n49__i1__net3 n63__i1__net3 125e-3
rk5627 n181__i1__i13__net1 n182__i1__i13__net1 75.287
rk5628 n182__i1__i13__net1 n183__i1__i13__net1 75.22e-3
rk5629 n183__i1__i13__net1 n184__i1__i13__net1 346e-3
rk5630 n181__i1__i13__net1 n183__i1__i13__net1 3.75
rk5632 n186__i1__i13__net1 n188__i1__i13__net1 186.7e-3
rk5633 n188__i1__i13__net1 n189__i1__i13__net1 151.2e-3
rk5634 n189__i1__i13__net1 n190__i1__i13__net1 323.1e-3
rk5635 n190__i1__i13__net1 n191__i1__i13__net1 57.75e-3
rk5636 n187__i1__i13__net1 n188__i1__i13__net1 3.1
rk5637 n187__i1__i13__net1 n191__i1__i13__net1 5.1667
rk5638 n51__i1__net3 n64__i1__net3 125e-3
rk5639 n53__i1__net3 n65__i1__net3 125e-3
rk5640 n1651__vss n1652__vss 115.8e-3
rk5641 n1652__vss n1653__vss 246.5e-3
rk5642 n1653__vss n1654__vss 97.36e-3
rk5644 n1651__vss n1656__vss 175.2e-3
rk5645 n1650__vss n1651__vss 75
rk5646 n1650__vss n1653__vss 3.75
rk5647 n1813__vddio n1814__vddio 459.3e-3
rk5648 n1814__vddio n1816__vddio 25.11e-3
rk5649 n1816__vddio n1817__vddio 318.7e-3
rk5650 n1817__vddio n1818__vddio 228e-3
rk5651 n1818__vddio n1819__vddio 190.3e-3
rk5652 n1815__vddio n1816__vddio 3.1
rk5653 n1815__vddio n1818__vddio 5.1667
rk5654 n1631__vddio n1820__vddio 2.5315
rk5655 n1820__vddio n1821__vddio 75.81e-3
rk5656 n1821__vddio n1822__vddio 73.24e-3
rk5657 n1822__vddio n1823__vddio 47.09e-3
rk5658 n1823__vddio n1824__vddio 145.3e-3
rk5659 n1824__vddio n1825__vddio 23.13e-3
rk5660 n1825__vddio n1826__vddio 290e-3
rk5661 n1826__vddio n1631__vddio 1.2852
rk5662 n1631__vddio n1821__vddio 1.25
rk5663 n1631__vddio n1823__vddio 1.25
rk5664 n1631__vddio n1825__vddio 1.25
rk5665 n1013__vss n1657__vss 2.0982
rk5666 n1657__vss n1658__vss 75.81e-3
rk5667 n1658__vss n1659__vss 73.24e-3
rk5668 n1659__vss n1660__vss 47.09e-3
rk5669 n1660__vss n1661__vss 145.3e-3
rk5670 n1661__vss n1662__vss 23.13e-3
rk5671 n1662__vss n1663__vss 290e-3
rk5672 n1663__vss n1013__vss 1.0686
rk5673 n1013__vss n1658__vss 1.0333
rk5674 n1013__vss n1660__vss 1.0333
rk5675 n1013__vss n1662__vss 1.0333
rl1 i1__i14__net1 n2__i1__i14__net1 22.9087
rl2 n3__i1__i14__net1 n4__i1__i14__net1 23.2215
rl3 n5__i1__i14__net1 n6__i1__i14__net1 22.8664
rl4 n7__i1__i14__net1 n8__i1__i14__net1 22.8664
rl5 n9__i1__i14__net1 n10__i1__i14__net1 23.2215
rl6 n11__i1__i14__net1 n12__i1__i14__net1 23.2215
rl7 n13__i1__i14__net1 n14__i1__i14__net1 22.8664
rl8 n15__i1__i14__net1 n16__i1__i14__net1 22.8664
rl9 n17__i1__i14__net1 n18__i1__i14__net1 23.2215
rl10 n19__i1__i14__net1 n20__i1__i14__net1 23.2215
rl11 i5__clk4 n2__i5__clk4 113.308
rl12 n2__i5__clk4 n3__i5__clk4 47.923
rl13 n4__i5__clk4 n5__i5__clk4 113.308
rl14 n5__i5__clk4 n6__i5__clk4 47.923
rl15 n21__i1__i14__net1 n22__i1__i14__net1 24.4918
rl16 n23__i1__i14__net1 n24__i1__i14__net1 24.4918
rl17 n25__i1__i14__net1 n26__i1__i14__net1 23.6861
rl18 n27__i1__i14__net1 n28__i1__i14__net1 23.6861
rl19 n1__x0 n2__x0 77.7258
rl20 n2__x0 n3__x0 45
rl21 n2__x0 n4__x0 104.649
rl22 n1__y0 n2__y0 77.7258
rl23 n2__y0 n3__y0 45
rl24 n2__y0 n4__y0 104.649
rl25 n29__i1__i14__net1 n30__i1__i14__net1 24.4918
rl26 n31__i1__i14__net1 n32__i1__i14__net1 24.4918
rl27 n33__i1__i14__net1 n34__i1__i14__net1 23.6861
rl28 n35__i1__i14__net1 n36__i1__i14__net1 23.6861
rl29 n7__i5__clk4 n8__i5__clk4 86.0764
rl30 i5__i7__i0__net1 n2__i5__i7__i0__net1 87.9995
rl31 n9__i5__clk4 n10__i5__clk4 86.0764
rl32 i5__i7__i1__net1 n2__i5__i7__i1__net1 87.9995
rl33 n37__i1__i14__net1 n38__i1__i14__net1 24.4918
rl34 n39__i1__i14__net1 n40__i1__i14__net1 24.4918
rl35 n41__i1__i14__net1 n42__i1__i14__net1 23.6861
rl36 n43__i1__i14__net1 n44__i1__i14__net1 23.6861
rl37 i5__i7__i0__i3__net22 n2__i5__i7__i0__i3__net22 77.7258
rl38 n2__i5__i7__i0__i3__net22 n3__i5__i7__i0__i3__net22 45
rl39 n2__i5__i7__i0__i3__net22 n4__i5__i7__i0__i3__net22 104.649
rl40 i5__i7__i1__i3__net22 n2__i5__i7__i1__i3__net22 77.7258
rl41 n2__i5__i7__i1__i3__net22 n3__i5__i7__i1__i3__net22 45
rl42 n2__i5__i7__i1__i3__net22 n4__i5__i7__i1__i3__net22 104.649
rl43 n45__i1__i14__net1 n46__i1__i14__net1 24.4918
rl44 n47__i1__i14__net1 n48__i1__i14__net1 24.4918
rl45 n3__i5__i7__i0__net1 n4__i5__i7__i0__net1 86.0764
rl46 n11__i5__clk4 n12__i5__clk4 87.9995
rl47 n3__i5__i7__i1__net1 n4__i5__i7__i1__net1 86.0764
rl48 n13__i5__clk4 n14__i5__clk4 87.9995
rl49 n49__i1__i14__net1 n50__i1__i14__net1 23.6861
rl50 n51__i1__i14__net1 n52__i1__i14__net1 23.6861
rl51 n53__i1__i14__net1 n54__i1__i14__net1 24.4918
rl52 n55__i1__i14__net1 n56__i1__i14__net1 24.4918
rl53 n1__reset n2__reset 82.2302
rl54 n3__reset n4__reset 82.2302
rl55 n57__i1__i14__net1 n58__i1__i14__net1 23.6861
rl56 n59__i1__i14__net1 n60__i1__i14__net1 23.6861
rl57 n65__i1__i14__net1 n66__i1__i14__net1 24.4918
rl58 n67__i1__i14__net1 n68__i1__i14__net1 24.4918
rl59 n1__x1 n2__x1 77.7258
rl60 n2__x1 n3__x1 45
rl61 n2__x1 n4__x1 104.649
rl62 n1__y1 n2__y1 77.7258
rl63 n2__y1 n3__y1 45
rl64 n2__y1 n4__y1 104.649
rl65 n77__i1__i14__net1 n78__i1__i14__net1 23.6861
rl66 n79__i1__i14__net1 n80__i1__i14__net1 23.6861
rl67 n15__i5__clk4 n16__i5__clk4 86.0764
rl68 n5__i5__i7__i0__net1 n6__i5__i7__i0__net1 87.9995
rl69 n81__i1__i14__net1 n82__i1__i14__net1 23.2215
rl70 n83__i1__i14__net1 n84__i1__i14__net1 23.2215
rl71 n17__i5__clk4 n18__i5__clk4 86.0764
rl72 n5__i5__i7__i1__net1 n6__i5__i7__i1__net1 87.9995
rl73 n89__i1__i14__net1 n90__i1__i14__net1 23.6861
rl74 n91__i1__i14__net1 n92__i1__i14__net1 23.6861
rl75 i5__i7__i0__i0__net22 n2__i5__i7__i0__i0__net22 77.7258
rl76 n2__i5__i7__i0__i0__net22 n3__i5__i7__i0__i0__net22 45
rl77 n2__i5__i7__i0__i0__net22 n4__i5__i7__i0__i0__net22 104.649
rl78 i5__i7__i1__i0__net22 n2__i5__i7__i1__i0__net22 77.7258
rl79 n2__i5__i7__i1__i0__net22 n3__i5__i7__i1__i0__net22 45
rl80 n2__i5__i7__i1__i0__net22 n4__i5__i7__i1__i0__net22 104.649
rl81 n97__i1__i14__net1 n98__i1__i14__net1 23.2215
rl82 n99__i1__i14__net1 n100__i1__i14__net1 23.2215
rl83 n105__i1__i14__net1 n106__i1__i14__net1 23.6861
rl84 n107__i1__i14__net1 n108__i1__i14__net1 23.6861
rl85 n11__i5__i7__i0__net1 n12__i5__i7__i0__net1 86.0764
rl86 n26__i5__clk4 n27__i5__clk4 87.9995
rl87 n11__i5__i7__i1__net1 n12__i5__i7__i1__net1 86.0764
rl88 n28__i5__clk4 n29__i5__clk4 87.9995
rl89 n113__i1__i14__net1 n114__i1__i14__net1 23.2215
rl90 n115__i1__i14__net1 n116__i1__i14__net1 23.2215
rl91 n125__i1__i14__net1 n126__i1__i14__net1 23.6861
rl92 n127__i1__i14__net1 n128__i1__i14__net1 23.6861
rl93 n5__reset n6__reset 82.2302
rl94 n7__reset n8__reset 82.2302
rl95 n131__i1__i14__net1 n132__i1__i14__net1 23.2215
rl96 n133__i1__i14__net1 n134__i1__i14__net1 23.2215
rl97 n1__x2 n2__x2 77.7258
rl98 n2__x2 n3__x2 45
rl99 n2__x2 n4__x2 104.649
rl100 n1__y2 n2__y2 77.7258
rl101 n2__y2 n3__y2 45
rl102 n2__y2 n4__y2 104.649
rl103 n141__i1__i14__net1 n142__i1__i14__net1 23.6861
rl104 n143__i1__i14__net1 n144__i1__i14__net1 23.6861
rl105 n145__i1__i14__net1 n146__i1__i14__net1 23.2215
rl106 n147__i1__i14__net1 n148__i1__i14__net1 23.2215
rl107 n36__i5__clk4 n37__i5__clk4 86.0764
rl108 n16__i5__i7__i0__net1 n17__i5__i7__i0__net1 87.9995
rl109 n38__i5__clk4 n39__i5__clk4 86.0764
rl110 n16__i5__i7__i1__net1 n17__i5__i7__i1__net1 87.9995
rl111 n157__i1__i14__net1 n158__i1__i14__net1 23.6861
rl112 n159__i1__i14__net1 n160__i1__i14__net1 23.6861
rl113 n161__i1__i14__net1 n162__i1__i14__net1 23.2215
rl114 n163__i1__i14__net1 n164__i1__i14__net1 23.2215
rl115 i5__i7__i0__i1__net22 n2__i5__i7__i0__i1__net22 77.7258
rl116 n2__i5__i7__i0__i1__net22 n3__i5__i7__i0__i1__net22 45
rl117 n2__i5__i7__i0__i1__net22 n4__i5__i7__i0__i1__net22 104.649
rl118 i5__i7__i1__i1__net22 n2__i5__i7__i1__i1__net22 77.7258
rl119 n2__i5__i7__i1__i1__net22 n3__i5__i7__i1__i1__net22 45
rl120 n2__i5__i7__i1__i1__net22 n4__i5__i7__i1__i1__net22 104.649
rl121 n173__i1__i14__net1 n174__i1__i14__net1 23.6861
rl122 n175__i1__i14__net1 n176__i1__i14__net1 23.6861
rl123 n18__i5__i7__i0__net1 n19__i5__i7__i0__net1 86.0764
rl124 n40__i5__clk4 n41__i5__clk4 87.9995
rl125 n18__i5__i7__i1__net1 n19__i5__i7__i1__net1 86.0764
rl126 n42__i5__clk4 n43__i5__clk4 87.9995
rl127 n177__i1__i14__net1 n178__i1__i14__net1 23.2215
rl128 n179__i1__i14__net1 n180__i1__i14__net1 23.2215
rl129 n185__i1__i14__net1 n186__i1__i14__net1 23.6861
rl130 n187__i1__i14__net1 n188__i1__i14__net1 23.6861
rl131 n16__reset n17__reset 82.2302
rl132 n18__reset n19__reset 82.2302
rl133 n197__i1__i14__net1 n198__i1__i14__net1 23.2215
rl134 n199__i1__i14__net1 n200__i1__i14__net1 23.2215
rl135 n201__i1__i14__net1 n202__i1__i14__net1 23.6861
rl136 n203__i1__i14__net1 n204__i1__i14__net1 23.6861
rl137 n1__x3 n2__x3 77.7258
rl138 n2__x3 n3__x3 45
rl139 n2__x3 n4__x3 104.649
rl140 n1__y3 n2__y3 77.7258
rl141 n2__y3 n3__y3 45
rl142 n2__y3 n4__y3 104.649
rl143 n209__i1__i14__net1 n210__i1__i14__net1 23.2215
rl144 n211__i1__i14__net1 n212__i1__i14__net1 23.2215
rl145 n217__i1__i14__net1 n218__i1__i14__net1 23.2215
rl146 n219__i1__i14__net1 n220__i1__i14__net1 23.2215
rl147 n46__i5__clk4 n47__i5__clk4 86.0764
rl148 n21__i5__i7__i0__net1 n22__i5__i7__i0__net1 87.9995
rl149 n48__i5__clk4 n49__i5__clk4 86.0764
rl150 n21__i5__i7__i1__net1 n22__i5__i7__i1__net1 87.9995
rl151 n225__i1__i14__net1 n226__i1__i14__net1 23.2215
rl152 n227__i1__i14__net1 n228__i1__i14__net1 23.2215
rl153 i5__i7__i0__i2__net22 n2__i5__i7__i0__i2__net22 77.7258
rl154 n2__i5__i7__i0__i2__net22 n3__i5__i7__i0__i2__net22 45
rl155 n2__i5__i7__i0__i2__net22 n4__i5__i7__i0__i2__net22 104.649
rl156 i5__i7__i1__i2__net22 n2__i5__i7__i1__i2__net22 77.7258
rl157 n2__i5__i7__i1__i2__net22 n3__i5__i7__i1__i2__net22 45
rl158 n2__i5__i7__i1__i2__net22 n4__i5__i7__i1__i2__net22 104.649
rl159 n237__i1__i14__net1 n238__i1__i14__net1 23.2215
rl160 n239__i1__i14__net1 n240__i1__i14__net1 23.2215
rl161 n241__i1__i14__net1 n242__i1__i14__net1 23.2215
rl162 n243__i1__i14__net1 n244__i1__i14__net1 23.2215
rl163 n25__i5__i7__i0__net1 n26__i5__i7__i0__net1 86.0764
rl164 n54__i5__clk4 n55__i5__clk4 87.9995
rl165 n25__i5__i7__i1__net1 n26__i5__i7__i1__net1 86.0764
rl166 n56__i5__clk4 n57__i5__clk4 87.9995
rl167 n253__i1__i14__net1 n254__i1__i14__net1 23.2215
rl168 n255__i1__i14__net1 n256__i1__i14__net1 23.2215
rl169 n257__i1__i14__net1 n258__i1__i14__net1 23.2215
rl170 n259__i1__i14__net1 n260__i1__i14__net1 23.2215
rl171 n24__reset n25__reset 82.2302
rl172 n26__reset n27__reset 82.2302
rl173 n269__i1__i14__net1 n270__i1__i14__net1 23.2215
rl174 n271__i1__i14__net1 n272__i1__i14__net1 23.2215
rl175 n273__i1__i14__net1 n274__i1__i14__net1 23.2215
rl176 n275__i1__i14__net1 n276__i1__i14__net1 23.2215
rl177 i5__i7__y2out n2__i5__i7__y2out 113.308
rl178 n2__i5__i7__y2out n3__i5__i7__y2out 47.923
rl179 n8__i5__i7__y1out n9__i5__i7__y1out 113.308
rl180 n9__i5__i7__y1out n10__i5__i7__y1out 47.923
rl181 n285__i1__i14__net1 n286__i1__i14__net1 23.6861
rl182 n287__i1__i14__net1 n288__i1__i14__net1 23.6861
rl183 n293__i1__i14__net1 n294__i1__i14__net1 23.2215
rl184 n295__i1__i14__net1 n296__i1__i14__net1 23.2215
rl185 i5__i7__x2out n2__i5__i7__x2out 80.7692
rl186 n2__i5__i7__x2out n3__i5__i7__x2out 103.022
rl187 n8__i5__i7__x1out n9__i5__i7__x1out 80.7692
rl188 n9__i5__i7__x1out n10__i5__i7__x1out 103.022
rl189 n301__i1__i14__net1 n302__i1__i14__net1 23.6861
rl190 n303__i1__i14__net1 n304__i1__i14__net1 23.6861
rl191 n305__i1__i14__net1 n306__i1__i14__net1 24.4918
rl192 n307__i1__i14__net1 n308__i1__i14__net1 24.4918
rl193 n11__i5__i7__y2out n12__i5__i7__y2out 66.6736
rl194 i5__i7__i8__net1 n2__i5__i7__i8__net1 108.981
rl195 n11__i5__i7__y1out n12__i5__i7__y1out 66.6736
rl196 i5__i7__i3__net1 n2__i5__i7__i3__net1 108.981
rl197 n313__i1__i14__net1 n314__i1__i14__net1 23.6861
rl198 n315__i1__i14__net1 n316__i1__i14__net1 23.6861
rl199 n325__i1__i14__net1 n326__i1__i14__net1 24.4918
rl200 n327__i1__i14__net1 n328__i1__i14__net1 24.4918
rl201 n333__i1__i14__net1 n334__i1__i14__net1 23.6861
rl202 n335__i1__i14__net1 n336__i1__i14__net1 23.6861
rl203 i5__i7__y3out n2__i5__i7__y3out 113.308
rl204 n2__i5__i7__y3out n3__i5__i7__y3out 47.923
rl205 n8__i5__i7__y0out n9__i5__i7__y0out 113.308
rl206 n9__i5__i7__y0out n10__i5__i7__y0out 47.923
rl207 n341__i1__i14__net1 n342__i1__i14__net1 24.4918
rl208 n343__i1__i14__net1 n344__i1__i14__net1 24.4918
rl209 n345__i1__i14__net1 n346__i1__i14__net1 23.6861
rl210 n347__i1__i14__net1 n348__i1__i14__net1 23.6861
rl211 i5__i7__x3out n2__i5__i7__x3out 80.7692
rl212 n2__i5__i7__x3out n3__i5__i7__x3out 103.022
rl213 n8__i5__i7__x0out n9__i5__i7__x0out 80.7692
rl214 n9__i5__i7__x0out n10__i5__i7__x0out 103.022
rl215 n357__i1__i14__net1 n358__i1__i14__net1 24.4918
rl216 n359__i1__i14__net1 n360__i1__i14__net1 24.4918
rl217 n361__i1__i14__net1 n362__i1__i14__net1 23.6861
rl218 n363__i1__i14__net1 n364__i1__i14__net1 23.6861
rl219 n4__i5__i7__y3out n5__i5__i7__y3out 66.6736
rl220 i5__i7__i9__net1 n2__i5__i7__i9__net1 108.981
rl221 n11__i5__i7__y0out n12__i5__i7__y0out 66.6736
rl222 i5__i7__i2__net1 n2__i5__i7__i2__net1 108.981
rl223 n373__i1__i14__net1 n374__i1__i14__net1 24.4918
rl224 n375__i1__i14__net1 n376__i1__i14__net1 24.4918
rl225 n379__i1__i14__net1 n380__i1__i14__net1 23.6861
rl226 n381__i1__i14__net1 n382__i1__i14__net1 23.6861
rl227 n389__i1__i14__net1 n390__i1__i14__net1 24.4918
rl228 n391__i1__i14__net1 n392__i1__i14__net1 24.4918
rl229 i5__i7__xor2 n2__i5__i7__xor2 113.308
rl230 n2__i5__i7__xor2 n3__i5__i7__xor2 47.923
rl231 i5__i7__xor1 n2__i5__i7__xor1 113.308
rl232 n2__i5__i7__xor1 n3__i5__i7__xor1 47.923
rl233 n393__i1__i14__net1 n394__i1__i14__net1 23.6861
rl234 n395__i1__i14__net1 n396__i1__i14__net1 23.6861
rl235 n405__i1__i14__net1 n406__i1__i14__net1 24.4918
rl236 n407__i1__i14__net1 n408__i1__i14__net1 24.4918
rl237 n413__i1__i14__net1 n414__i1__i14__net1 23.6861
rl238 n415__i1__i14__net1 n416__i1__i14__net1 23.6861
rl239 i5__i7__i5__net1 n2__i5__i7__i5__net1 86.0245
rl240 n2__i5__i7__i5__net1 n3__i5__i7__i5__net1 11.25
rl241 n2__i5__i7__i5__net1 n4__i5__i7__i5__net1 112.948
rl242 i5__i7__i4__net1 n2__i5__i7__i4__net1 86.0245
rl243 n2__i5__i7__i4__net1 n3__i5__i7__i4__net1 11.25
rl244 n2__i5__i7__i4__net1 n4__i5__i7__i4__net1 112.948
rl245 n421__i1__i14__net1 n422__i1__i14__net1 24.4918
rl246 n423__i1__i14__net1 n424__i1__i14__net1 24.4918
rl247 n425__i1__i14__net1 n426__i1__i14__net1 23.6861
rl248 n427__i1__i14__net1 n428__i1__i14__net1 23.6861
rl249 n11__i5__i7__xor2 n12__i5__i7__xor2 102.04
rl250 n11__i5__i7__xor1 n12__i5__i7__xor1 102.04
rl251 n433__i1__i14__net1 n434__i1__i14__net1 23.2215
rl252 n435__i1__i14__net1 n436__i1__i14__net1 23.2215
rl253 n441__i1__i14__net1 n442__i1__i14__net1 23.6861
rl254 n443__i1__i14__net1 n444__i1__i14__net1 23.6861
rl255 i5__i7__xor3 n2__i5__i7__xor3 80.7692
rl256 n2__i5__i7__xor3 n3__i5__i7__xor3 103.022
rl257 i5__i7__xor0 n2__i5__i7__xor0 80.7692
rl258 n2__i5__i7__xor0 n3__i5__i7__xor0 103.022
rl259 n449__i1__i14__net1 n450__i1__i14__net1 23.2215
rl260 n451__i1__i14__net1 n452__i1__i14__net1 23.2215
rl261 n457__i1__i14__net1 n458__i1__i14__net1 23.6861
rl262 n459__i1__i14__net1 n460__i1__i14__net1 23.6861
rl263 n13__i5__i7__xor2 n14__i5__i7__xor2 66.6736
rl264 n5__i5__i7__i5__net1 n6__i5__i7__i5__net1 108.981
rl265 n13__i5__i7__xor1 n14__i5__i7__xor1 66.6736
rl266 n5__i5__i7__i4__net1 n6__i5__i7__i4__net1 108.981
rl267 n465__i1__i14__net1 n466__i1__i14__net1 23.2215
rl268 n467__i1__i14__net1 n468__i1__i14__net1 23.2215
rl269 n477__i1__i14__net1 n478__i1__i14__net1 23.6861
rl270 n479__i1__i14__net1 n480__i1__i14__net1 23.6861
rl271 n481__i1__i14__net1 n482__i1__i14__net1 23.2215
rl272 n483__i1__i14__net1 n484__i1__i14__net1 23.2215
rl273 i5__i7__net51 n2__i5__i7__net51 113.308
rl274 n2__i5__i7__net51 n3__i5__i7__net51 47.923
rl275 i5__i7__net47 n2__i5__i7__net47 113.308
rl276 n2__i5__i7__net47 n3__i5__i7__net47 47.923
rl277 n493__i1__i14__net1 n494__i1__i14__net1 23.6861
rl278 n495__i1__i14__net1 n496__i1__i14__net1 23.6861
rl279 n497__i1__i14__net1 n498__i1__i14__net1 23.2215
rl280 n499__i1__i14__net1 n500__i1__i14__net1 23.2215
rl281 i5__i7__net44 n2__i5__i7__net44 80.7692
rl282 n2__i5__i7__net44 n3__i5__i7__net44 103.022
rl283 n505__i1__i14__net1 n506__i1__i14__net1 23.6861
rl284 n507__i1__i14__net1 n508__i1__i14__net1 23.6861
rl285 i5__i7__i6__net1 n2__i5__i7__i6__net1 86.0245
rl286 n2__i5__i7__i6__net1 n3__i5__i7__i6__net1 11.25
rl287 n2__i5__i7__i6__net1 n4__i5__i7__i6__net1 112.948
rl288 n513__i1__i14__net1 n514__i1__i14__net1 23.2215
rl289 n515__i1__i14__net1 n516__i1__i14__net1 23.2215
rl290 n4__i5__i7__net47 n5__i5__i7__net47 66.6736
rl291 i5__i7__i7__i0__net1 n2__i5__i7__i7__i0__net1 108.981
rl292 n525__i1__i14__net1 n526__i1__i14__net1 23.6861
rl293 n527__i1__i14__net1 n528__i1__i14__net1 23.6861
rl294 n4__i5__i7__net51 n5__i5__i7__net51 102.04
rl295 n529__i1__i14__net1 n530__i1__i14__net1 23.2215
rl296 n531__i1__i14__net1 n532__i1__i14__net1 23.2215
rl297 i5__i7__net50 n2__i5__i7__net50 80.7692
rl298 n2__i5__i7__net50 n3__i5__i7__net50 103.022
rl299 n541__i1__i14__net1 n542__i1__i14__net1 23.2215
rl300 n543__i1__i14__net1 n544__i1__i14__net1 23.2215
rl301 i5__i7__i7__net1 n2__i5__i7__i7__net1 113.308
rl302 n2__i5__i7__i7__net1 n3__i5__i7__i7__net1 47.923
rl303 n545__i1__i14__net1 n546__i1__i14__net1 23.2215
rl304 n547__i1__i14__net1 n548__i1__i14__net1 23.2215
rl305 n6__i5__i7__net51 n7__i5__i7__net51 66.6736
rl306 n5__i5__i7__i6__net1 n6__i5__i7__i6__net1 108.981
rl307 n553__i1__i14__net1 n554__i1__i14__net1 23.2215
rl308 n555__i1__i14__net1 n556__i1__i14__net1 23.2215
rl309 n561__i1__i14__net1 n562__i1__i14__net1 23.2215
rl310 n563__i1__i14__net1 n564__i1__i14__net1 23.2215
rl311 i5__i7__net46 n2__i5__i7__net46 80.7692
rl312 n2__i5__i7__net46 n3__i5__i7__net46 103.022
rl313 n569__i1__i14__net1 n570__i1__i14__net1 23.2215
rl314 n571__i1__i14__net1 n572__i1__i14__net1 23.2215
rl315 i5__clk_buf n2__i5__clk_buf 88.4156
rl316 n2__i5__clk_buf n3__i5__clk_buf 88.5818
rl317 n3__i5__clk_buf n4__i5__clk_buf 82.2455
rl318 n2__i5__clk_buf n5__i5__clk_buf 21.372
rl319 n4__i5__clk_buf n6__i5__clk_buf 82.2455
rl320 n6__i5__clk_buf n7__i5__clk_buf 88.4156
rl321 n7__i5__clk_buf n8__i5__clk_buf 21.372
rl322 n7__i5__clk_buf n9__i5__clk_buf 88.5818
rl323 n577__i1__i14__net1 n578__i1__i14__net1 23.2215
rl324 n579__i1__i14__net1 n580__i1__i14__net1 23.2215
rl325 n4__i5__i7__i7__net1 n5__i5__i7__i7__net1 66.6736
rl326 i5__i7__i7__i1__net1 n2__i5__i7__i7__i1__net1 108.981
rl327 n589__i1__i14__net1 n590__i1__i14__net1 23.2215
rl328 n591__i1__i14__net1 n592__i1__i14__net1 23.2215
rl329 n1__shift n2__shift 49.8461
rl330 n2__shift n3__shift 88.3077
rl331 n593__i1__i14__net1 n594__i1__i14__net1 23.2215
rl332 n595__i1__i14__net1 n596__i1__i14__net1 23.2215
rl333 n6__i5__i7__i7__net1 n7__i5__i7__i7__net1 113.308
rl334 n7__i5__i7__i7__net1 n8__i5__i7__i7__net1 47.923
rl335 n605__i1__i14__net1 n606__i1__i14__net1 23.2215
rl336 n607__i1__i14__net1 n608__i1__i14__net1 23.2215
rl337 i5__i6__i6__net4 n2__i5__i6__i6__net4 80.3072
rl338 n4__shift n5__shift 89.9225
rl339 n609__i1__i14__net1 n610__i1__i14__net1 23.2215
rl340 n611__i1__i14__net1 n612__i1__i14__net1 23.2215
rl341 n617__i1__i14__net1 n618__i1__i14__net1 23.2215
rl342 n619__i1__i14__net1 n620__i1__i14__net1 23.2215
rl343 n6__shift n7__shift 89.9225
rl344 n3__i5__i6__i6__net4 n4__i5__i6__i6__net4 80.3072
rl345 i5__i7__i7__net2 n2__i5__i7__i7__net2 71.5013
rl346 n10__i5__i7__net44 n11__i5__i7__net44 71.5013
rl347 n629__i1__i14__net1 n630__i1__i14__net1 23.2215
rl348 n631__i1__i14__net1 n632__i1__i14__net1 23.2215
rl349 n637__i1__i14__net1 n638__i1__i14__net1 23.2215
rl350 n639__i1__i14__net1 n640__i1__i14__net1 23.2215
rl351 n8__i5__i7__net46 n9__i5__i7__net46 71.5013
rl352 n3__i5__i7__i7__net2 n4__i5__i7__i7__net2 71.5013
rl353 i5__i6__net30 n2__i5__i6__net30 83.1872
rl354 n2__i5__i6__net30 n3__i5__i6__net30 43.2071
rl355 n3__i5__i6__net30 n4__i5__i6__net30 39.3609
rl356 n4__i5__i6__net30 n5__i5__i6__net30 26.8981
rl357 n2__i5__i6__net30 n6__i5__i6__net30 26.8981
rl358 n4__i5__i6__net30 n7__i5__i6__net30 83.3534
rl359 n645__i1__i14__net1 n646__i1__i14__net1 23.2215
rl360 n647__i1__i14__net1 n648__i1__i14__net1 23.2215
rl361 n14__i5__i7__i7__net1 n15__i5__i7__i7__net1 73.9763
rl362 n10__i5__i7__net46 n11__i5__i7__net46 67.6551
rl363 n10__i5__clk_buf n11__i5__clk_buf 109.826
rl364 n11__i5__clk_buf n12__i5__clk_buf 86.5405
rl365 i5__i6__net31 n2__i5__i6__net31 81.3628
rl366 n2__i5__i6__net31 n3__i5__i6__net31 55.5169
rl367 n2__i5__i6__net31 n4__i5__i6__net31 26.3061
rl368 n649__i1__i14__net1 n650__i1__i14__net1 23.2215
rl369 n651__i1__i14__net1 n652__i1__i14__net1 23.2215
rl370 n19__i5__i7__net44 n20__i5__i7__net44 73.9763
rl371 n17__i5__i7__i7__net1 n18__i5__i7__i7__net1 73.9763
rl372 n657__i1__i14__net1 n658__i1__i14__net1 23.6861
rl373 n659__i1__i14__net1 n660__i1__i14__net1 23.6861
rl374 n669__i1__i14__net1 n670__i1__i14__net1 23.2215
rl375 n671__i1__i14__net1 n672__i1__i14__net1 23.2215
rl376 i5__i6__i2__net22 n2__i5__i6__i2__net22 83.1872
rl377 n2__i5__i6__i2__net22 n3__i5__i6__i2__net22 43.2071
rl378 n3__i5__i6__i2__net22 n4__i5__i6__i2__net22 39.3609
rl379 n4__i5__i6__i2__net22 n5__i5__i6__i2__net22 26.8981
rl380 n2__i5__i6__i2__net22 n6__i5__i6__i2__net22 26.8981
rl381 n4__i5__i6__i2__net22 n7__i5__i6__i2__net22 83.3534
rl382 n673__i1__i14__net1 n674__i1__i14__net1 23.6861
rl383 n675__i1__i14__net1 n676__i1__i14__net1 23.6861
rl384 i5__i7__i7__net3 n2__i5__i7__i7__net3 113.308
rl385 n2__i5__i7__i7__net3 n3__i5__i7__i7__net3 47.923
rl386 n5__i5__i6__net31 n6__i5__i6__net31 109.826
rl387 n6__i5__i6__net31 n7__i5__i6__net31 86.5405
rl388 n13__i5__clk_buf n14__i5__clk_buf 109.826
rl389 n14__i5__clk_buf n15__i5__clk_buf 86.5405
rl390 n685__i1__i14__net1 n686__i1__i14__net1 23.2215
rl391 n687__i1__i14__net1 n688__i1__i14__net1 23.2215
rl392 n689__i1__i14__net1 n690__i1__i14__net1 23.6861
rl393 n691__i1__i14__net1 n692__i1__i14__net1 23.6861
rl394 n36__reset n37__reset 96.7685
rl395 n37__reset n38__reset 111.662
rl396 n37__reset n39__reset 23.5864
rl397 n1__clk_out n2__clk_out 178.846
rl398 n2__clk_out n3__clk_out 109.826
rl399 n3__clk_out n4__clk_out 77.6148
rl400 n4__clk_out n5__clk_out 75.6918
rl401 n5__clk_out n6__clk_out 108.732
rl402 n6__clk_out n1__clk_out 9.1667
rl403 n701__i1__i14__net1 n702__i1__i14__net1 23.2215
rl404 n703__i1__i14__net1 n704__i1__i14__net1 23.2215
rl405 n705__i1__i14__net1 n706__i1__i14__net1 23.6861
rl406 n707__i1__i14__net1 n708__i1__i14__net1 23.6861
rl407 n10__shift n11__shift 49.8461
rl408 n11__shift n12__shift 88.3077
rl409 i5__i9__net21 n2__i5__i9__net21 82.2302
rl410 n2__i5__i9__net21 n3__i5__i9__net21 46.8456
rl411 n3__i5__i9__net21 n4__i5__i9__net21 46.8456
rl412 n4__i5__i9__net21 n5__i5__i9__net21 80.3072
rl413 n713__i1__i14__net1 n714__i1__i14__net1 23.2215
rl414 n715__i1__i14__net1 n716__i1__i14__net1 23.2215
rl415 n6__i5__i9__net21 n7__i5__i9__net21 82.2302
rl416 n8__i5__i9__net21 n9__i5__i9__net21 80.3072
rl417 n10__i5__i9__net21 n11__i5__i9__net21 82.2302
rl418 n12__i5__i9__net21 n13__i5__i9__net21 80.3072
rl419 i5__i6__i7__net4 n2__i5__i6__i7__net4 80.3072
rl420 n17__shift n18__shift 89.9225
rl421 n14__i5__i9__net21 n15__i5__i9__net21 82.2302
rl422 n16__i5__i9__net21 n17__i5__i9__net21 80.3072
rl423 n19__shift n20__shift 89.9225
rl424 n3__i5__i6__i7__net4 n4__i5__i6__i7__net4 80.3072
rl425 n18__i5__clk_buf n19__i5__clk_buf 88.4156
rl426 n19__i5__clk_buf n20__i5__clk_buf 88.5818
rl427 n20__i5__clk_buf n21__i5__clk_buf 82.2455
rl428 n19__i5__clk_buf n22__i5__clk_buf 21.372
rl429 n21__i5__clk_buf n23__i5__clk_buf 82.2455
rl430 n23__i5__clk_buf n24__i5__clk_buf 88.4156
rl431 n24__i5__clk_buf n25__i5__clk_buf 21.372
rl432 n24__i5__clk_buf n26__i5__clk_buf 88.5818
rl433 i5__i6__net33 n2__i5__i6__net33 83.1872
rl434 n2__i5__i6__net33 n3__i5__i6__net33 43.2071
rl435 n3__i5__i6__net33 n4__i5__i6__net33 39.3609
rl436 n4__i5__i6__net33 n5__i5__i6__net33 26.8981
rl437 n2__i5__i6__net33 n6__i5__i6__net33 26.8981
rl438 n4__i5__i6__net33 n7__i5__i6__net33 83.3534
rl439 n29__i5__clk_buf n30__i5__clk_buf 109.826
rl440 n30__i5__clk_buf n31__i5__clk_buf 86.5405
rl441 n18__i5__i6__net31 n19__i5__i6__net31 81.3628
rl442 n19__i5__i6__net31 n20__i5__i6__net31 55.5169
rl443 n19__i5__i6__net31 n21__i5__i6__net31 26.3061
rl444 i5__i8__net1 n2__i5__i8__net1 83.1872
rl445 n2__i5__i8__net1 n3__i5__i8__net1 43.2071
rl446 n3__i5__i8__net1 n4__i5__i8__net1 39.3609
rl447 n4__i5__i8__net1 n5__i5__i8__net1 26.8981
rl448 n2__i5__i8__net1 n6__i5__i8__net1 26.8981
rl449 n4__i5__i8__net1 n7__i5__i8__net1 83.3534
rl450 i1__net2 n2__i1__net2 24.4918
rl451 n3__i1__net2 n4__i1__net2 24.4918
rl452 n32__i5__clk_buf n33__i5__clk_buf 109.826
rl453 n33__i5__clk_buf n34__i5__clk_buf 86.5405
rl454 i5__i8__net4 n2__i5__i8__net4 81.3628
rl455 n2__i5__i8__net4 n3__i5__i8__net4 55.5169
rl456 n2__i5__i8__net4 n4__i5__i8__net4 26.3061
rl457 i5__i6__i4__net22 n2__i5__i6__i4__net22 83.1872
rl458 n2__i5__i6__i4__net22 n3__i5__i6__i4__net22 43.2071
rl459 n3__i5__i6__i4__net22 n4__i5__i6__i4__net22 39.3609
rl460 n4__i5__i6__i4__net22 n5__i5__i6__i4__net22 26.8981
rl461 n2__i5__i6__i4__net22 n6__i5__i6__i4__net22 26.8981
rl462 n4__i5__i6__i4__net22 n7__i5__i6__i4__net22 83.3534
rl463 n5__i1__net2 n6__i1__net2 23.6861
rl464 n7__i1__net2 n8__i1__net2 23.6861
rl465 n26__i5__i6__net31 n27__i5__i6__net31 109.826
rl466 n27__i5__i6__net31 n28__i5__i6__net31 86.5405
rl467 n37__i5__clk_buf n38__i5__clk_buf 109.826
rl468 n38__i5__clk_buf n39__i5__clk_buf 86.5405
rl469 n9__i1__net2 n10__i1__net2 24.4918
rl470 n11__i1__net2 n12__i1__net2 24.4918
rl471 i5__i8__i9__net22 n2__i5__i8__i9__net22 83.1872
rl472 n2__i5__i8__i9__net22 n3__i5__i8__i9__net22 43.2071
rl473 n3__i5__i8__i9__net22 n4__i5__i8__i9__net22 39.3609
rl474 n4__i5__i8__i9__net22 n5__i5__i8__i9__net22 26.8981
rl475 n2__i5__i8__i9__net22 n6__i5__i8__i9__net22 26.8981
rl476 n4__i5__i8__i9__net22 n7__i5__i8__i9__net22 83.3534
rl477 n13__i1__net2 n14__i1__net2 23.6861
rl478 n15__i1__net2 n16__i1__net2 23.6861
rl479 n5__i5__i8__net4 n6__i5__i8__net4 109.826
rl480 n6__i5__i8__net4 n7__i5__i8__net4 86.5405
rl481 n40__i5__clk_buf n41__i5__clk_buf 109.826
rl482 n41__i5__clk_buf n42__i5__clk_buf 86.5405
rl483 n17__i1__net2 n18__i1__net2 23.2215
rl484 n19__i1__net2 n20__i1__net2 23.2215
rl485 n43__reset n44__reset 96.7685
rl486 n44__reset n45__reset 111.662
rl487 n44__reset n46__reset 23.5864
rl488 n21__i1__net2 n22__i1__net2 23.6861
rl489 n23__i1__net2 n24__i1__net2 23.6861
rl490 n25__i1__net2 n26__i1__net2 23.2215
rl491 n27__i1__net2 n28__i1__net2 23.2215
rl492 n23__shift n24__shift 49.8461
rl493 n24__shift n25__shift 88.3077
rl494 n47__reset n48__reset 96.7685
rl495 n48__reset n49__reset 111.662
rl496 n48__reset n50__reset 23.5864
rl497 n29__i1__net2 n30__i1__net2 23.6861
rl498 n31__i1__net2 n32__i1__net2 23.6861
rl499 i5__i6__i8__net4 n2__i5__i6__i8__net4 80.3072
rl500 n30__shift n31__shift 89.9225
rl501 n33__i1__net2 n34__i1__net2 23.2215
rl502 n35__i1__net2 n36__i1__net2 23.2215
rl503 n37__i1__net2 n38__i1__net2 23.6861
rl504 n39__i1__net2 n40__i1__net2 23.6861
rl505 i5__i8__net2 n2__i5__i8__net2 88.4156
rl506 n2__i5__i8__net2 n3__i5__i8__net2 88.5818
rl507 n3__i5__i8__net2 n4__i5__i8__net2 82.2455
rl508 n2__i5__i8__net2 n5__i5__i8__net2 21.372
rl509 n4__i5__i8__net2 n6__i5__i8__net2 82.2455
rl510 n6__i5__i8__net2 n7__i5__i8__net2 88.4156
rl511 n7__i5__i8__net2 n8__i5__i8__net2 21.372
rl512 n7__i5__i8__net2 n9__i5__i8__net2 88.5818
rl513 n32__shift n33__shift 89.9225
rl514 n3__i5__i6__i8__net4 n4__i5__i6__i8__net4 80.3072
rl515 n41__i1__net2 n42__i1__net2 23.2215
rl516 n43__i1__net2 n44__i1__net2 23.2215
rl517 n45__i1__net2 n46__i1__net2 23.6861
rl518 n47__i1__net2 n48__i1__net2 23.6861
rl519 i5__i6__net35 n2__i5__i6__net35 83.1872
rl520 n2__i5__i6__net35 n3__i5__i6__net35 43.2071
rl521 n3__i5__i6__net35 n4__i5__i6__net35 39.3609
rl522 n4__i5__i6__net35 n5__i5__i6__net35 26.8981
rl523 n2__i5__i6__net35 n6__i5__i6__net35 26.8981
rl524 n4__i5__i6__net35 n7__i5__i6__net35 83.3534
rl525 i5__i8__net5 n2__i5__i8__net5 83.1872
rl526 n2__i5__i8__net5 n3__i5__i8__net5 43.2071
rl527 n3__i5__i8__net5 n4__i5__i8__net5 39.3609
rl528 n4__i5__i8__net5 n5__i5__i8__net5 26.8981
rl529 n2__i5__i8__net5 n6__i5__i8__net5 26.8981
rl530 n4__i5__i8__net5 n7__i5__i8__net5 83.3534
rl531 n49__i1__net2 n50__i1__net2 23.2215
rl532 n51__i1__net2 n52__i1__net2 23.2215
rl533 n53__i5__clk_buf n54__i5__clk_buf 109.826
rl534 n54__i5__clk_buf n55__i5__clk_buf 86.5405
rl535 n32__i5__i6__net31 n33__i5__i6__net31 81.3628
rl536 n33__i5__i6__net31 n34__i5__i6__net31 55.5169
rl537 n33__i5__i6__net31 n35__i5__i6__net31 26.3061
rl538 n53__i1__net2 n54__i1__net2 23.6861
rl539 n55__i1__net2 n56__i1__net2 23.6861
rl540 n10__i5__i8__net2 n11__i5__i8__net2 109.826
rl541 n11__i5__i8__net2 n12__i5__i8__net2 86.5405
rl542 n11__i5__i8__net1 n12__i5__i8__net1 81.3628
rl543 n12__i5__i8__net1 n13__i5__i8__net1 55.5169
rl544 n12__i5__i8__net1 n14__i5__i8__net1 26.3061
rl545 n57__i1__net2 n58__i1__net2 23.2215
rl546 n59__i1__net2 n60__i1__net2 23.2215
rl547 n65__i1__net2 n66__i1__net2 23.6861
rl548 n67__i1__net2 n68__i1__net2 23.6861
rl549 i5__i6__i5__net22 n2__i5__i6__i5__net22 83.1872
rl550 n2__i5__i6__i5__net22 n3__i5__i6__i5__net22 43.2071
rl551 n3__i5__i6__i5__net22 n4__i5__i6__i5__net22 39.3609
rl552 n4__i5__i6__i5__net22 n5__i5__i6__i5__net22 26.8981
rl553 n2__i5__i6__i5__net22 n6__i5__i6__i5__net22 26.8981
rl554 n4__i5__i6__i5__net22 n7__i5__i6__i5__net22 83.3534
rl555 i5__i8__i10__net22 n2__i5__i8__i10__net22 83.1872
rl556 n2__i5__i8__i10__net22 n3__i5__i8__i10__net22 43.2071
rl557 n3__i5__i8__i10__net22 n4__i5__i8__i10__net22 39.3609
rl558 n4__i5__i8__i10__net22 n5__i5__i8__i10__net22 26.8981
rl559 n2__i5__i8__i10__net22 n6__i5__i8__i10__net22 26.8981
rl560 n4__i5__i8__i10__net22 n7__i5__i8__i10__net22 83.3534
rl561 n73__i1__net2 n74__i1__net2 23.2215
rl562 n75__i1__net2 n76__i1__net2 23.2215
rl563 n38__i5__i6__net31 n39__i5__i6__net31 109.826
rl564 n39__i5__i6__net31 n40__i5__i6__net31 86.5405
rl565 n60__i5__clk_buf n61__i5__clk_buf 109.826
rl566 n61__i5__clk_buf n62__i5__clk_buf 86.5405
rl567 n15__i5__i8__net1 n16__i5__i8__net1 109.826
rl568 n16__i5__i8__net1 n17__i5__i8__net1 86.5405
rl569 n13__i5__i8__net2 n14__i5__i8__net2 109.826
rl570 n14__i5__i8__net2 n15__i5__i8__net2 86.5405
rl571 n85__i1__net2 n86__i1__net2 23.6861
rl572 n87__i1__net2 n88__i1__net2 23.6861
rl573 n93__i1__net2 n94__i1__net2 23.2215
rl574 n95__i1__net2 n96__i1__net2 23.2215
rl575 n56__reset n57__reset 96.7685
rl576 n57__reset n58__reset 111.662
rl577 n57__reset n59__reset 23.5864
rl578 n60__reset n61__reset 96.7685
rl579 n61__reset n62__reset 111.662
rl580 n61__reset n63__reset 23.5864
rl581 n101__i1__net2 n102__i1__net2 23.6861
rl582 n103__i1__net2 n104__i1__net2 23.6861
rl583 n105__i1__net2 n106__i1__net2 23.2215
rl584 n107__i1__net2 n108__i1__net2 23.2215
rl585 bufin n2__bufin 76.4763
rl586 n2__bufin n3__bufin 72.6302
rl587 n113__i1__net2 n114__i1__net2 23.2215
rl588 n115__i1__net2 n116__i1__net2 23.2215
rl589 n76__i5__clk4 n77__i5__clk4 88.4156
rl590 n77__i5__clk4 n78__i5__clk4 88.5818
rl591 n78__i5__clk4 n79__i5__clk4 82.2455
rl592 n77__i5__clk4 n80__i5__clk4 21.372
rl593 n79__i5__clk4 n81__i5__clk4 82.2455
rl594 n81__i5__clk4 n82__i5__clk4 88.4156
rl595 n82__i5__clk4 n83__i5__clk4 21.372
rl596 n82__i5__clk4 n84__i5__clk4 88.5818
rl597 n121__i1__net2 n122__i1__net2 23.2215
rl598 n123__i1__net2 n124__i1__net2 23.2215
rl599 i4__net1 n2__i4__net1 178.846
rl600 n2__i4__net1 n3__i4__net1 109.826
rl601 n3__i4__net1 n4__i4__net1 77.6148
rl602 n4__i4__net1 n5__i4__net1 75.6918
rl603 n5__i4__net1 n6__i4__net1 108.732
rl604 n6__i4__net1 i4__net1 9.1667
rl605 n133__i1__net2 n134__i1__net2 23.2215
rl606 n135__i1__net2 n136__i1__net2 23.2215
rl607 n85__i5__clk4 n86__i5__clk4 75.8027
rl608 n86__i5__clk4 n87__i5__clk4 46.8551
rl609 n86__i5__clk4 n88__i5__clk4 70.0334
rl610 n137__i1__net2 n138__i1__net2 23.2215
rl611 n139__i1__net2 n140__i1__net2 23.2215
rl612 n30__i5__i8__net2 n31__i5__i8__net2 155.769
rl613 n31__i5__i8__net2 n32__i5__i8__net2 98.4704
rl614 n145__i1__net2 n146__i1__net2 23.2215
rl615 n147__i1__net2 n148__i1__net2 23.2215
rl616 n1__piso_out n2__piso_out 110.772
rl617 n2__piso_out n3__piso_out 68.5478
rl618 n3__piso_out n4__piso_out 72.348
rl619 n4__piso_out n5__piso_out 75.7689
rl620 n5__piso_out n6__piso_out 13.7551
rl621 n2__piso_out n7__piso_out 118.464
rl622 n3__piso_out n8__piso_out 116.943
rl623 n3__piso_out n9__piso_out 109.251
rl624 n4__piso_out n10__piso_out 116.943
rl625 n4__piso_out n11__piso_out 109.251
rl626 n5__piso_out n12__piso_out 106.191
rl627 n5__piso_out n13__piso_out 104.268
rl628 n153__i1__net2 n154__i1__net2 23.2215
rl629 n155__i1__net2 n156__i1__net2 23.2215
rl630 i5__i8__i8__net1 n2__i5__i8__i8__net1 59.4615
rl631 n2__i5__i8__i8__net1 n3__i5__i8__i8__net1 46
rl632 n181__i1__net2 n182__i1__net2 23.2215
rl633 n183__i1__net2 n184__i1__net2 23.2215
rl634 i1__i13__net1 n2__i1__i13__net1 23.2215
rl635 n3__i1__i13__net1 n4__i1__i13__net1 23.2215
rl636 i1__i12__net1 n2__i1__i12__net1 23.6861
rl637 n3__i1__i12__net1 n4__i1__i12__net1 23.6861
rl638 n5__i1__i13__net1 n6__i1__i13__net1 23.2215
rl639 n7__i1__i13__net1 n8__i1__i13__net1 23.6861
rl640 n5__i1__i12__net1 n6__i1__i12__net1 23.6861
rl641 n7__i1__i12__net1 n8__i1__i12__net1 23.6861
rl642 n9__i1__i13__net1 n10__i1__i13__net1 23.2215
rl643 n11__i1__i13__net1 n12__i1__i13__net1 23.2215
rl644 n9__i1__i12__net1 n10__i1__i12__net1 23.6861
rl645 n11__i1__i12__net1 n12__i1__i12__net1 23.6861
rl646 n13__i1__i13__net1 n14__i1__i13__net1 23.2215
rl647 n15__i1__i13__net1 n16__i1__i13__net1 23.6861
rl648 n13__i1__i12__net1 n14__i1__i12__net1 23.6861
rl649 n15__i1__i12__net1 n16__i1__i12__net1 23.6861
rl650 n17__i1__i13__net1 n18__i1__i13__net1 23.2215
rl651 n19__i1__i13__net1 n20__i1__i13__net1 23.2215
rl652 n17__i1__i12__net1 n18__i1__i12__net1 23.6861
rl653 n19__i1__i12__net1 n20__i1__i12__net1 23.6861
rl654 n21__i1__i13__net1 n22__i1__i13__net1 23.6861
rl655 n23__i1__i13__net1 n24__i1__i13__net1 23.6861
rl656 n21__i1__i12__net1 n22__i1__i12__net1 23.6861
rl657 n23__i1__i12__net1 n24__i1__i12__net1 23.6861
rl658 n25__i1__i13__net1 n26__i1__i13__net1 23.2215
rl659 n27__i1__i13__net1 n28__i1__i13__net1 24.4918
rl660 n25__i1__i12__net1 n26__i1__i12__net1 23.6861
rl661 n27__i1__i12__net1 n28__i1__i12__net1 23.6861
rl662 n29__i1__i13__net1 n30__i1__i13__net1 23.6861
rl663 n31__i1__i13__net1 n32__i1__i13__net1 23.6861
rl664 n33__i1__i13__net1 n34__i1__i13__net1 23.2215
rl665 n35__i1__i13__net1 n36__i1__i13__net1 24.4918
rl666 n37__i1__i13__net1 n38__i1__i13__net1 23.6861
rl667 n39__i1__i13__net1 n40__i1__i13__net1 23.6861
rl668 i1__net4 n2__i1__net4 23.6861
rl669 n3__i1__net4 n4__i1__net4 23.6861
rl670 n41__i1__i13__net1 n42__i1__i13__net1 23.2215
rl671 n43__i1__i13__net1 n44__i1__i13__net1 24.4918
rl672 n5__i1__net4 n6__i1__net4 23.6861
rl673 n7__i1__net4 n8__i1__net4 23.6861
rl674 n45__i1__i13__net1 n46__i1__i13__net1 23.6861
rl675 n47__i1__i13__net1 n48__i1__i13__net1 23.6861
rl676 n49__i1__i13__net1 n50__i1__i13__net1 23.2215
rl677 n51__i1__i13__net1 n52__i1__i13__net1 24.4918
rl678 n53__i1__i13__net1 n54__i1__i13__net1 23.6861
rl679 n55__i1__i13__net1 n56__i1__i13__net1 23.6861
rl681 n20__piso_out n22__piso_out 12.45
rl682 n20__piso_out n23__piso_out 26.3213
rl683 n9__i1__net4 n10__i1__net4 38.963
rl684 n57__i1__i13__net1 n58__i1__i13__net1 23.2215
rl685 n59__i1__i13__net1 n60__i1__i13__net1 24.4918
rl686 n24__piso_out n25__piso_out 38.963
rl687 n11__i1__net4 n12__i1__net4 38.963
rl688 n65__i1__i13__net1 n66__i1__i13__net1 23.6861
rl689 n67__i1__i13__net1 n68__i1__i13__net1 23.6861
rl690 n26__piso_out n27__piso_out 38.963
rl691 n77__i1__i13__net1 n78__i1__i13__net1 23.2215
rl692 n79__i1__i13__net1 n80__i1__i13__net1 24.4918
rl693 n81__i1__i13__net1 n82__i1__i13__net1 23.6861
rl694 n83__i1__i13__net1 n84__i1__i13__net1 23.6861
rl695 n9__piso_outinv n10__piso_outinv 37.0036
rl696 n89__i1__i13__net1 n90__i1__i13__net1 23.2215
rl697 n91__i1__i13__net1 n92__i1__i13__net1 24.4918
rl698 i1__i11__outinv n2__i1__i11__outinv 39.7609
rl699 n11__piso_outinv n12__piso_outinv 39.7609
rl700 n97__i1__i13__net1 n98__i1__i13__net1 23.6861
rl701 n99__i1__i13__net1 n100__i1__i13__net1 23.6861
rl702 n3__i1__i11__outinv n4__i1__i11__outinv 38.963
rl703 n13__piso_outinv n14__piso_outinv 39.7609
rl704 n121__i1__i13__net1 n122__i1__i13__net1 23.2215
rl705 n123__i1__i13__net1 n124__i1__i13__net1 24.4918
rl706 n30__i1__net3 n31__i1__net3 23.6861
rl707 n32__i1__net3 n33__i1__net3 23.6861
rl708 n34__i1__net3 n35__i1__net3 23.6861
rl709 n36__i1__net3 n37__i1__net3 23.6861
rl710 n38__i1__net3 n39__i1__net3 23.2215
rl711 n40__i1__net3 n41__i1__net3 23.2215
rl712 n42__i1__net3 n43__i1__net3 23.6861
rl713 n44__i1__net3 n45__i1__net3 23.6861
rl714 n46__i1__net3 n47__i1__net3 23.2215
rl715 n48__i1__net3 n49__i1__net3 23.2215
rl716 n50__i1__net3 n51__i1__net3 23.6861
rl717 n52__i1__net3 n53__i1__net3 23.6861
mi1__i14__m1_96__rcx n45__vddio n24__i1__i14__net1 n119__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_95__rcx n80__chipdriverout n19__i1__i14__net1 n45__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_94__rcx n24__vddio n15__i1__i14__net1 n80__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_93__rcx n41__chipdriverout n11__i1__i14__net1 n24__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_92__rcx n3__vddio n7__i1__i14__net1 n41__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_91__rcx n3__chipdriverout n3__i1__i14__net1 n3__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.44e-12 AS=1.44e-12 PD=19.55e-6 PS=19.55e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_90__rcx n118__vddio n48__i1__i14__net1 n247__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_89__rcx n208__chipdriverout n43__i1__i14__net1 n118__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_88__rcx n97__vddio n40__i1__i14__net1 n208__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_87__rcx n169__chipdriverout n35__i1__i14__net1 n97__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_86__rcx n70__vddio n32__i1__i14__net1 n169__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_85__rcx n119__chipdriverout n27__i1__i14__net1 n70__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_84__rcx n181__vddio n83__i1__i14__net1 n364__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_83__rcx n325__chipdriverout n79__i1__i14__net1 n181__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_82__rcx n160__vddio n68__i1__i14__net1 n325__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_81__rcx n286__chipdriverout n59__i1__i14__net1 n160__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_80__rcx n139__vddio n56__i1__i14__net1 n286__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_79__rcx n247__chipdriverout n51__i1__i14__net1 n139__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_78__rcx n254__vddio n133__i1__i14__net1 n470__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_77__rcx n442__chipdriverout n127__i1__i14__net1 n254__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_76__rcx n246__vddio n115__i1__i14__net1 n442__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_75__rcx n403__chipdriverout n107__i1__i14__net1 n246__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_74__rcx n212__vddio n99__i1__i14__net1 n403__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_73__rcx n364__chipdriverout n91__i1__i14__net1 n212__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_72__rcx n327__vddio n179__i1__i14__net1 n587__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_71__rcx n573__chipdriverout n175__i1__i14__net1 n327__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_70__rcx n319__vddio n163__i1__i14__net1 n573__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_69__rcx n534__chipdriverout n159__i1__i14__net1 n319__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_68__rcx n285__vddio n147__i1__i14__net1 n534__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_67__rcx n470__chipdriverout n143__i1__i14__net1 n285__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_66__rcx n403__vddio n227__i1__i14__net1 n704__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_65__rcx n665__chipdriverout n219__i1__i14__net1 n403__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_64__rcx n382__vddio n211__i1__i14__net1 n665__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_63__rcx n626__chipdriverout n203__i1__i14__net1 n382__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_62__rcx n361__vddio n199__i1__i14__net1 n626__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_61__rcx n587__chipdriverout n187__i1__i14__net1 n361__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_60__rcx n463__vddio n275__i1__i14__net1 n832__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_59__rcx n793__chipdriverout n271__i1__i14__net1 n463__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_58__rcx n449__vddio n259__i1__i14__net1 n793__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_57__rcx n743__chipdriverout n255__i1__i14__net1 n449__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_56__rcx n428__vddio n243__i1__i14__net1 n743__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_55__rcx n704__chipdriverout n239__i1__i14__net1 n428__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_54__rcx n526__vddio n328__i1__i14__net1 n949__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_53__rcx n910__chipdriverout n315__i1__i14__net1 n526__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_52__rcx n505__vddio n308__i1__i14__net1 n910__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_51__rcx n860__chipdriverout n303__i1__i14__net1 n505__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_50__rcx n484__vddio n295__i1__i14__net1 n860__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_49__rcx n832__chipdriverout n287__i1__i14__net1 n484__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_48__rcx n949__chipdriverout n335__i1__i14__net1 n560__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_47__rcx n1066__chipdriverout n381__i1__i14__net1 n620__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_46__rcx n612__vddio n376__i1__i14__net1 n1066__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_45__rcx n1027__chipdriverout n363__i1__i14__net1 n612__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_44__rcx n578__vddio n360__i1__i14__net1 n1027__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_43__rcx n1008__chipdriverout n347__i1__i14__net1 n578__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_42__rcx n560__vddio n344__i1__i14__net1 n1008__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_41__rcx n1183__chipdriverout n427__i1__i14__net1 n693__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_40__rcx n685__vddio n424__i1__i14__net1 n1183__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_39__rcx n1144__chipdriverout n415__i1__i14__net1 n685__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_38__rcx n651__vddio n408__i1__i14__net1 n1144__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_37__rcx n1125__chipdriverout n395__i1__i14__net1 n651__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_36__rcx n620__vddio n392__i1__i14__net1 n1125__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_35__rcx n1300__chipdriverout n479__i1__i14__net1 n756__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_34__rcx n735__vddio n467__i1__i14__net1 n1300__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_33__rcx n1261__chipdriverout n459__i1__i14__net1 n735__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_32__rcx n714__vddio n451__i1__i14__net1 n1261__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_31__rcx n1222__chipdriverout n443__i1__i14__net1 n714__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_30__rcx n693__vddio n435__i1__i14__net1 n1222__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_29__rcx n1417__chipdriverout n527__i1__i14__net1 n842__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_28__rcx n802__vddio n515__i1__i14__net1 n1417__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_27__rcx n1378__chipdriverout n507__i1__i14__net1 n802__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_26__rcx n777__vddio n499__i1__i14__net1 n1378__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_25__rcx n1339__chipdriverout n495__i1__i14__net1 n777__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_24__rcx n756__vddio n483__i1__i14__net1 n1339__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_23__rcx n1551__chipdriverout n571__i1__i14__net1 n892__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_22__rcx n884__vddio n563__i1__i14__net1 n1551__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_21__rcx n1511__chipdriverout n555__i1__i14__net1 n884__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_20__rcx n850__vddio n547__i1__i14__net1 n1511__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_19__rcx n1478__chipdriverout n543__i1__i14__net1 n850__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_18__rcx n842__vddio n531__i1__i14__net1 n1478__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_17__rcx n1658__chipdriverout n619__i1__i14__net1 n965__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_16__rcx n944__vddio n611__i1__i14__net1 n1658__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_15__rcx n1619__chipdriverout n607__i1__i14__net1 n944__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_14__rcx n923__vddio n595__i1__i14__net1 n1619__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_13__rcx n1591__chipdriverout n591__i1__i14__net1 n923__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_12__rcx n892__vddio n579__i1__i14__net1 n1591__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_11__rcx n1775__chipdriverout n671__i1__i14__net1 n1038__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_10__rcx n1020__vddio n659__i1__i14__net1 n1775__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_9__rcx n1736__chipdriverout n651__i1__i14__net1 n1020__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_8__rcx n986__vddio n647__i1__i14__net1 n1736__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_7__rcx n1697__chipdriverout n639__i1__i14__net1 n986__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_6__rcx n965__vddio n631__i1__i14__net1 n1697__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_5__rcx n1080__vddio n707__i1__i14__net1 n1892__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_4__rcx n1853__chipdriverout n703__i1__i14__net1 n1080__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_3__rcx n1059__vddio n691__i1__i14__net1 n1853__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_2__rcx n1830__chipdriverout n687__i1__i14__net1 n1059__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1_1__rcx n1038__vddio n675__i1__i14__net1 n1830__chipdriverout n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m1 n1892__chipdriverout n715__i1__i14__net1 n1101__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.55e-6 PS=19.55e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_27__rcx n1257__vddio n27__i1__net2 n921__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_26__rcx n882__i1__i14__net1 n23__i1__net2 n1257__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_25__rcx n1223__vddio n19__i1__net2 n882__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_24__rcx n843__i1__i14__net1 n15__i1__net2 n1223__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_23__rcx n1202__vddio n12__i1__net2 n843__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_22__rcx n804__i1__i14__net1 n7__i1__net2 n1202__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_21__rcx n1175__vddio n4__i1__net2 n804__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.44e-12 AS=1.44e-12 PD=19.55e-6 PS=19.55e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_20__rcx n1027__i1__i14__net1 n55__i1__net2 n1351__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_19__rcx n1317__vddio n51__i1__net2 n1027__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_18__rcx n999__i1__i14__net1 n47__i1__net2 n1317__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_17__rcx n1296__vddio n43__i1__net2 n999__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_16__rcx n960__i1__i14__net1 n39__i1__net2 n1296__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_15__rcx n1265__vddio n35__i1__net2 n960__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_14__rcx n921__i1__i14__net1 n31__i1__net2 n1265__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_13__rcx n1411__vddio n107__i1__net2 n1183__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_12__rcx n1155__i1__i14__net1 n103__i1__net2 n1411__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_11__rcx n1380__vddio n95__i1__net2 n1155__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_10__rcx n1116__i1__i14__net1 n87__i1__net2 n1380__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_9__rcx n1359__vddio n75__i1__net2 n1116__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_8__rcx n1091__i1__i14__net1 n67__i1__net2 n1359__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_7__rcx n1351__vddio n59__i1__net2 n1091__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_6__rcx n1331__i1__i14__net1 n183__i1__net2 n1523__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.55e-6 PS=19.55e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_5__rcx n1487__vddio n155__i1__net2 n1331__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_4__rcx n1272__i1__i14__net1 n147__i1__net2 n1487__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_3__rcx n1453__vddio n139__i1__net2 n1272__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_2__rcx n1222__i1__i14__net1 n135__i1__net2 n1453__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0_1__rcx n1432__vddio n123__i1__net2 n1222__i1__i14__net1 n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m0 n1183__i1__i14__net1 n115__i1__net2 n1432__vddio n1631__vddio g45p2svt L=150e-9 W=9.6e-6 AD=1.92e-12 AS=1.92e-12 PD=19.6e-6 PS=19.6e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i11__m2_1__rcx n8__i1__i11__outinv n12__i1__net4 n1784__vddio n1767__vddio g45p2svt L=150e-9 W=320e-9 AD=64e-15 AS=64e-15 PD=990e-9 PS=990e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i11__m2 n1778__vddio n10__i1__net4 n8__i1__i11__outinv n1767__vddio g45p2svt L=150e-9 W=320e-9 AD=48e-15 AS=48e-15 PD=990e-9 PS=990e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i11__m3_1__rcx n1776__vddio n2__i1__i11__outinv n26__i1__net4 n1767__vddio g45p2svt L=150e-9 W=320e-9 AD=48e-15 AS=48e-15 PD=990e-9 PS=990e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i11__m3 n26__i1__net4 n4__i1__i11__outinv n1766__vddio n1767__vddio g45p2svt L=150e-9 W=320e-9 AD=64e-15 AS=64e-15 PD=990e-9 PS=990e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_20__rcx n259__i1__net2 n25__i1__i13__net1 n1700__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_19__rcx n1693__vddio n21__i1__i13__net1 n259__i1__net2 n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_18__rcx n250__i1__net2 n17__i1__i13__net1 n1693__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_17__rcx n1686__vddio n13__i1__i13__net1 n250__i1__net2 n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_16__rcx n245__i1__net2 n9__i1__i13__net1 n1686__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_15__rcx n1679__vddio n5__i1__i13__net1 n245__i1__net2 n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_14__rcx n232__i1__net2 i1__i13__net1 n1679__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=576e-15 AS=576e-15 PD=8.03e-6 PS=8.03e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_13__rcx n1700__vddio n29__i1__i13__net1 n268__i1__net2 n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_12__rcx n295__i1__net2 n57__i1__i13__net1 n1746__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_11__rcx n1739__vddio n53__i1__i13__net1 n295__i1__net2 n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_10__rcx n286__i1__net2 n49__i1__i13__net1 n1739__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_9__rcx n1714__vddio n45__i1__i13__net1 n286__i1__net2 n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_8__rcx n277__i1__net2 n41__i1__i13__net1 n1714__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_7__rcx n1708__vddio n37__i1__i13__net1 n277__i1__net2 n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_6__rcx n268__i1__net2 n33__i1__i13__net1 n1708__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_5__rcx n326__i1__net2 n121__i1__i13__net1 n1786__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.03e-6 PS=8.03e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_4__rcx n1760__vddio n97__i1__i13__net1 n326__i1__net2 n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_3__rcx n317__i1__net2 n89__i1__i13__net1 n1760__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_2__rcx n1753__vddio n81__i1__i13__net1 n317__i1__net2 n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3_1__rcx n304__i1__net2 n77__i1__i13__net1 n1753__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m3 n1746__vddio n65__i1__i13__net1 n304__i1__net2 n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m2_5__rcx n187__i1__i13__net1 n52__i1__net3 n1815__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.03e-6 PS=8.03e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m2_4__rcx n1807__vddio n48__i1__net3 n187__i1__i13__net1 n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m2_3__rcx n176__i1__i13__net1 n44__i1__net3 n1807__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m2_2__rcx n1800__vddio n40__i1__net3 n176__i1__i13__net1 n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m2_1__rcx n165__i1__i13__net1 n36__i1__net3 n1800__vddio n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=768e-15 AS=768e-15 PD=8.08e-6 PS=8.08e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m2 n1794__vddio n32__i1__net3 n165__i1__i13__net1 n1631__vddio g45p2svt L=150e-9 W=3.84e-6 AD=576e-15 AS=576e-15 PD=8.03e-6 PS=8.03e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m1_1__rcx n62__i1__i12__net1 n7__i1__net4 n1779__vddio n1767__vddio g45p2svt L=150e-9 W=960e-9 AD=192e-15 AS=192e-15 PD=2.27e-6 PS=2.27e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m1 n1780__vddio n3__i1__net4 n62__i1__i12__net1 n1767__vddio g45p2svt L=150e-9 W=960e-9 AD=144e-15 AS=144e-15 PD=2.27e-6 PS=2.27e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m0_6__rcx n24__i1__net3 n27__i1__i12__net1 n1781__vddio n1767__vddio g45p2svt L=150e-9 W=960e-9 AD=192e-15 AS=192e-15 PD=2.27e-6 PS=2.27e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m0_5__rcx n1782__vddio n23__i1__i12__net1 n24__i1__net3 n1767__vddio g45p2svt L=150e-9 W=960e-9 AD=192e-15 AS=192e-15 PD=2.32e-6 PS=2.32e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m0_4__rcx n19__i1__net3 n19__i1__i12__net1 n1782__vddio n1767__vddio g45p2svt L=150e-9 W=960e-9 AD=192e-15 AS=192e-15 PD=2.32e-6 PS=2.32e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m0_3__rcx n1783__vddio n15__i1__i12__net1 n19__i1__net3 n1767__vddio g45p2svt L=150e-9 W=960e-9 AD=192e-15 AS=192e-15 PD=2.32e-6 PS=2.32e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m0_2__rcx n12__i1__net3 n11__i1__i12__net1 n1783__vddio n1767__vddio g45p2svt L=150e-9 W=960e-9 AD=192e-15 AS=192e-15 PD=2.32e-6 PS=2.32e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m0_1__rcx n1775__vddio n7__i1__i12__net1 n12__i1__net3 n1767__vddio g45p2svt L=150e-9 W=960e-9 AD=192e-15 AS=192e-15 PD=2.32e-6 PS=2.32e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m0 n4__i1__net3 n3__i1__i12__net1 n1775__vddio n1767__vddio g45p2svt L=150e-9 W=960e-9 AD=144e-15 AS=144e-15 PD=2.27e-6 PS=2.27e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi5__i8__i5__pm0_2__rcx n13__i5__i8__net5 n76__i5__clk4 n270__vdd n182__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i5__pm0_1__rcx n18__i5__i8__net5 n78__i5__clk4 n271__vdd n182__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i5__pm0 n270__vdd n80__i5__clk4 n18__i5__i8__net5 n182__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i4__pm0_2__rcx n18__i5__i8__net1 i5__i8__net2 n274__vdd n182__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i4__pm0_1__rcx n23__i5__i8__net1 n3__i5__i8__net2 n275__vdd n182__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i4__pm0 n274__vdd n5__i5__i8__net2 n23__i5__i8__net1 n182__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i6__pm0_2__rcx n8__i5__i8__net4 n18__i5__clk_buf n278__vdd n182__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i6__pm0_1__rcx n14__i5__i8__net4 n20__i5__clk_buf n279__vdd n182__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i6__pm0 n278__vdd n22__i5__clk_buf n14__i5__i8__net4 n182__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__pm1_1__rcx n272__vdd n6__i5__i8__i10__net22 i5__i8__i10__net24 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__pm1 n4__i5__i8__i10__net24 i5__i8__i10__net22 n272__vdd n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__pm0_1__rcx n97__i5__clk4 n16__i5__i8__net1 n4__i5__i8__i10__net24 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__pm0 n7__i5__i8__i10__net24 n15__i5__i8__net1 n97__i5__clk4 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__pm3_1__rcx n273__vdd n6__i5__i8__net5 i5__i8__i10__net25 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__pm3 n4__i5__i8__i10__net25 i5__i8__net5 n273__vdd n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__pm2_1__rcx n8__i5__i8__i10__net22 n11__i5__i8__net2 n4__i5__i8__i10__net25 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__pm2 n8__i5__i8__i10__net25 n10__i5__i8__net2 n8__i5__i8__i10__net22 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__pm1_1__rcx n276__vdd n6__i5__i8__i9__net22 i5__i8__i9__net24 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__pm1 n4__i5__i8__i9__net24 i5__i8__i9__net22 n276__vdd n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__pm0_1__rcx n29__i5__i8__net2 n6__i5__i8__net4 n4__i5__i8__i9__net24 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__pm0 n8__i5__i8__i9__net24 n5__i5__i8__net4 n29__i5__i8__net2 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__pm3_1__rcx n277__vdd n6__i5__i8__net1 i5__i8__i9__net25 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__pm3 n4__i5__i8__i9__net25 i5__i8__net1 n277__vdd n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__pm2_1__rcx n8__i5__i8__i9__net22 n33__i5__clk_buf n4__i5__i8__i9__net25 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__pm2 n7__i5__i8__i9__net25 n32__i5__clk_buf n8__i5__i8__i9__net22 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i8__pm2 n44__shift i5__i8__i8__net1 n181__vdd n182__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i8__pm0 i5__i8__i8__net2 n85__i5__clk4 n269__vdd n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i8__pm1 n4__i5__i8__i8__net1 n30__i5__i8__net2 i5__i8__i8__net2 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i2__pm1 n2__i5__i7__i1__i2__net24 i5__i7__i1__i2__net22 n291__vdd n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i2__pm0 n8__i5__i7__y3out n25__i5__i7__i1__net1 i5__i7__i1__i2__net24 n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i2__pm3 n2__i5__i7__i1__i2__net21 n1__y3 n292__vdd n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i2__pm2 n5__i5__i7__i1__i2__net22 n48__i5__clk4 i5__i7__i1__i2__net21 n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i1__pm1 n2__i5__i7__i1__i1__net24 i5__i7__i1__i1__net22 n293__vdd n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i1__pm0 n6__i5__i7__y2out n18__i5__i7__i1__net1 i5__i7__i1__i1__net24 n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i1__pm3 n2__i5__i7__i1__i1__net21 n1__y2 n294__vdd n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i1__pm2 n5__i5__i7__i1__i1__net22 n38__i5__clk4 i5__i7__i1__i1__net21 n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i0__pm1 n2__i5__i7__i1__i0__net24 i5__i7__i1__i0__net22 n295__vdd n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i0__pm0 n3__i5__i7__y1out n11__i5__i7__i1__net1 i5__i7__i1__i0__net24 n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i0__pm3 n2__i5__i7__i1__i0__net21 n1__y1 n296__vdd n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i0__pm2 n5__i5__i7__i1__i0__net22 n17__i5__clk4 i5__i7__i1__i0__net21 n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i3__pm1 n2__i5__i7__i1__i3__net24 i5__i7__i1__i3__net22 n297__vdd n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i3__pm0 n3__i5__i7__y0out n3__i5__i7__i1__net1 i5__i7__i1__i3__net24 n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i3__pm3 n2__i5__i7__i1__i3__net21 n1__y0 n298__vdd n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i3__pm2 n5__i5__i7__i1__i3__net22 n9__i5__clk4 i5__i7__i1__i3__net21 n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i4__pm0 n9__i5__i7__i1__net1 n4__i5__clk4 n299__vdd n237__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i2__pm1 n2__i5__i7__i0__i2__net24 i5__i7__i0__i2__net22 n308__vdd n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i2__pm0 n6__i5__i7__x3out n25__i5__i7__i0__net1 i5__i7__i0__i2__net24 n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i2__pm3 n2__i5__i7__i0__i2__net21 n1__x3 n307__vdd n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i2__pm2 n5__i5__i7__i0__i2__net22 n46__i5__clk4 i5__i7__i0__i2__net21 n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i1__pm1 n2__i5__i7__i0__i1__net24 i5__i7__i0__i1__net22 n306__vdd n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i1__pm0 n6__i5__i7__x2out n18__i5__i7__i0__net1 i5__i7__i0__i1__net24 n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i1__pm3 n2__i5__i7__i0__i1__net21 n1__x2 n305__vdd n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i1__pm2 n5__i5__i7__i0__i1__net22 n36__i5__clk4 i5__i7__i0__i1__net21 n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i0__pm1 n2__i5__i7__i0__i0__net24 i5__i7__i0__i0__net22 n304__vdd n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i0__pm0 n3__i5__i7__x1out n11__i5__i7__i0__net1 i5__i7__i0__i0__net24 n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i0__pm3 n2__i5__i7__i0__i0__net21 n1__x1 n303__vdd n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i0__pm2 n5__i5__i7__i0__i0__net22 n15__i5__clk4 i5__i7__i0__i0__net21 n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i3__pm1 n2__i5__i7__i0__i3__net24 i5__i7__i0__i3__net22 n302__vdd n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i3__pm0 n3__i5__i7__x0out n3__i5__i7__i0__net1 i5__i7__i0__i3__net24 n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i3__pm3 n2__i5__i7__i0__i3__net21 n1__x0 n301__vdd n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i3__pm2 n5__i5__i7__i0__i3__net22 n7__i5__clk4 i5__i7__i0__i3__net21 n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i4__pm0 n9__i5__i7__i0__net1 i5__clk4 n300__vdd n256__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i5__i0__pm0 n8__i5__i7__net47 i5__i7__i5__net1 n10__i5__i7__xor3 n221__vdd g45p1svt L=45e-9 W=240e-9 AD=46.8e-15 AS=46.8e-15 PD=875e-9 PS=875e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i5__i1__pm0 n23__i5__i7__xor3 n13__i5__i7__xor2 n8__i5__i7__net51 n221__vdd g45p1svt L=45e-9 W=240e-9 AD=54e-15 AS=54e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i5__i1__pm1 n8__i5__i7__net51 i5__i7__xor3 n22__i5__i7__xor2 n221__vdd g45p1svt L=45e-9 W=240e-9 AD=133.2e-15 AS=133.2e-15 PD=1.265e-6 PS=1.265e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i5__i2__pm0 n7__i5__i7__i5__net1 i5__i7__xor2 n288__vdd n221__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i6__i0__pm0 n6__i5__i7__net46 i5__i7__i6__net1 n10__i5__i7__net50 n328__vdd g45p1svt L=45e-9 W=240e-9 AD=46.8e-15 AS=46.8e-15 PD=875e-9 PS=875e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i6__i1__pm0 n21__i5__i7__net50 n6__i5__i7__net51 n4__i5__r0 n328__vdd g45p1svt L=45e-9 W=240e-9 AD=54e-15 AS=54e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i6__i1__pm1 n4__i5__r0 i5__i7__net50 n22__i5__i7__net51 n328__vdd g45p1svt L=45e-9 W=240e-9 AD=133.2e-15 AS=133.2e-15 PD=1.265e-6 PS=1.265e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i6__i2__pm0 n9__i5__i7__i6__net1 i5__i7__net51 n327__vdd n328__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i4__i0__pm0 n6__i5__i7__net44 i5__i7__i4__net1 n10__i5__i7__xor0 n322__vdd g45p1svt L=45e-9 W=240e-9 AD=46.8e-15 AS=46.8e-15 PD=875e-9 PS=875e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i4__i1__pm0 n23__i5__i7__xor0 n13__i5__i7__xor1 n4__i5__i7__net50 n322__vdd g45p1svt L=45e-9 W=240e-9 AD=54e-15 AS=54e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i4__i1__pm1 n4__i5__i7__net50 i5__i7__xor0 n22__i5__i7__xor1 n322__vdd g45p1svt L=45e-9 W=240e-9 AD=133.2e-15 AS=133.2e-15 PD=1.265e-6 PS=1.265e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i4__i2__pm0 n7__i5__i7__i4__net1 i5__i7__xor1 n321__vdd n322__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i1__i0__pm0 n14__i5__i7__net46 n4__i5__i7__i7__net1 i5__r1 n182__vdd g45p1svt L=45e-9 W=240e-9 AD=54e-15 AS=54e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i1__i0__pm1 i5__r1 i5__i7__net46 n20__i5__i7__i7__net1 n182__vdd g45p1svt L=45e-9 W=240e-9 AD=133.2e-15 AS=133.2e-15 PD=1.265e-6 PS=1.265e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i1__i1__pm0 n3__i5__i7__i7__i1__net1 i5__i7__i7__net1 n286__vdd n182__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i0__i0__pm0 n13__i5__i7__net44 n4__i5__i7__net47 n9__i5__i7__i7__net1 n182__vdd g45p1svt L=45e-9 W=240e-9 AD=54e-15 AS=54e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i0__i0__pm1 n9__i5__i7__i7__net1 i5__i7__net44 n13__i5__i7__net47 n182__vdd g45p1svt L=45e-9 W=240e-9 AD=133.2e-15 AS=133.2e-15 PD=1.265e-6 PS=1.265e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i0__i1__pm0 n3__i5__i7__i7__i0__net1 i5__i7__net47 n287__vdd n182__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i4__pm0 i5__i7__i7__i4__net2 i5__i7__i7__net2 n284__vdd n182__vdd g45p1svt L=45e-9 W=240e-9 AD=75.6e-15 AS=75.6e-15 PD=1.005e-6 PS=1.005e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i4__pm1 n4__i5__i7__i7__net3 n8__i5__i7__net46 i5__i7__i7__i4__net2 n182__vdd g45p1svt L=45e-9 W=240e-9 AD=75.6e-15 AS=75.6e-15 PD=1.11e-6 PS=1.11e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i4__pm3 i5__i7__i7__i4__net3 n15__i5__i7__i7__net1 n4__i5__i7__i7__net3 n182__vdd g45p1svt L=45e-9 W=240e-9 AD=75.6e-15 AS=75.6e-15 PD=1.11e-6 PS=1.11e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i4__pm2 n283__vdd n20__i5__i7__net44 i5__i7__i7__i4__net3 n182__vdd g45p1svt L=45e-9 W=240e-9 AD=54e-15 AS=54e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i2__pm0 n5__i5__i7__i7__net2 n6__i5__i7__i7__net1 n285__vdd n182__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i3__pm0 n10__i5__r2 i5__i7__i7__net3 n282__vdd n182__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i9__i0__pm0 n14__i5__i7__x3out n4__i5__i7__y3out n4__i5__i7__xor3 n228__vdd g45p1svt L=45e-9 W=240e-9 AD=54e-15 AS=54e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i9__i0__pm1 n4__i5__i7__xor3 i5__i7__x3out n15__i5__i7__y3out n228__vdd g45p1svt L=45e-9 W=240e-9 AD=133.2e-15 AS=133.2e-15 PD=1.265e-6 PS=1.265e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i9__i1__pm0 n3__i5__i7__i9__net1 i5__i7__y3out n289__vdd n228__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i8__i0__pm0 n14__i5__i7__x2out n11__i5__i7__y2out n4__i5__i7__xor2 n233__vdd g45p1svt L=45e-9 W=240e-9 AD=54e-15 AS=54e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i8__i0__pm1 n4__i5__i7__xor2 i5__i7__x2out n17__i5__i7__y2out n233__vdd g45p1svt L=45e-9 W=240e-9 AD=133.2e-15 AS=133.2e-15 PD=1.265e-6 PS=1.265e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i8__i1__pm0 n3__i5__i7__i8__net1 i5__i7__y2out n290__vdd n233__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i2__i0__pm0 n14__i5__i7__x0out n11__i5__i7__y0out n4__i5__i7__xor0 n317__vdd g45p1svt L=45e-9 W=240e-9 AD=54e-15 AS=54e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i2__i0__pm1 n4__i5__i7__xor0 n8__i5__i7__x0out n17__i5__i7__y0out n317__vdd g45p1svt L=45e-9 W=240e-9 AD=133.2e-15 AS=133.2e-15 PD=1.265e-6 PS=1.265e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i2__i1__pm0 n3__i5__i7__i2__net1 n8__i5__i7__y0out n316__vdd n317__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i3__i0__pm0 n14__i5__i7__x1out n11__i5__i7__y1out n4__i5__i7__xor1 n312__vdd g45p1svt L=45e-9 W=240e-9 AD=54e-15 AS=54e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i3__i0__pm1 n4__i5__i7__xor1 n8__i5__i7__x1out n17__i5__i7__y1out n312__vdd g45p1svt L=45e-9 W=240e-9 AD=133.2e-15 AS=133.2e-15 PD=1.265e-6 PS=1.265e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i3__i1__pm0 n3__i5__i7__i3__net1 n8__i5__i7__y1out n311__vdd n312__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i9__pm1_3__rcx n161__vdd n15__i5__i9__net21 n49__i5__clk_buf n182__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i9__pm0_1__rcx n18__i5__i9__net21 n5__clk_out n281__vdd n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i9__pm0 n280__vdd n1__clk_out n18__i5__i9__net21 n182__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i9__pm1_2__rcx n50__i5__clk_buf n2__i5__i9__net21 n152__vdd n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i9__pm1_1__rcx n155__vdd n7__i5__i9__net21 n50__i5__clk_buf n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i9__pm1 n49__i5__clk_buf n11__i5__i9__net21 n155__vdd n182__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i9__pm0_2__rcx n8__i5__i6__net31 i5__clk_buf n336__vdd n328__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i9__pm0_1__rcx n14__i5__i6__net31 n3__i5__clk_buf n333__vdd n328__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i9__pm0 n336__vdd n5__i5__clk_buf n14__i5__i6__net31 n328__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__pm1_1__rcx n362__vdd n6__i5__i6__i5__net22 i5__i6__i5__net24 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__pm1 n4__i5__i6__i5__net24 i5__i6__i5__net22 n362__vdd n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__pm0_1__rcx n10__bufin n39__i5__i6__net31 n4__i5__i6__i5__net24 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__pm0 n8__i5__i6__i5__net24 n38__i5__i6__net31 n10__bufin n328__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__pm3_1__rcx n359__vdd n6__i5__i6__net35 i5__i6__i5__net25 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__pm3 n4__i5__i6__i5__net25 i5__i6__net35 n359__vdd n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__pm2_1__rcx n8__i5__i6__i5__net22 n54__i5__clk_buf n4__i5__i6__i5__net25 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__pm2 n8__i5__i6__i5__net25 n53__i5__clk_buf n8__i5__i6__i5__net22 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__pm1_1__rcx n353__vdd n6__i5__i6__i4__net22 i5__i6__i4__net24 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__pm1 n4__i5__i6__i4__net24 i5__i6__i4__net22 n353__vdd n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__pm0_1__rcx n7__i5__i6__net34 n27__i5__i6__net31 n4__i5__i6__i4__net24 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__pm0 n7__i5__i6__i4__net24 n26__i5__i6__net31 n7__i5__i6__net34 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__pm3_1__rcx n350__vdd n6__i5__i6__net33 i5__i6__i4__net25 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__pm3 n4__i5__i6__i4__net25 i5__i6__net33 n350__vdd n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__pm2_1__rcx n8__i5__i6__i4__net22 n30__i5__clk_buf n4__i5__i6__i4__net25 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__pm2 n7__i5__i6__i4__net25 n29__i5__clk_buf n8__i5__i6__i4__net22 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__pm1_1__rcx n344__vdd n6__i5__i6__i2__net22 i5__i6__i2__net24 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__pm1 n4__i5__i6__i2__net24 i5__i6__i2__net22 n344__vdd n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__pm0_1__rcx n7__i5__i6__net32 n6__i5__i6__net31 n4__i5__i6__i2__net24 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__pm0 n7__i5__i6__i2__net24 n5__i5__i6__net31 n7__i5__i6__net32 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__pm3_1__rcx n341__vdd n6__i5__i6__net30 i5__i6__i2__net25 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__pm3 n4__i5__i6__i2__net25 i5__i6__net30 n341__vdd n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__pm2_1__rcx n8__i5__i6__i2__net22 n11__i5__clk_buf n4__i5__i6__i2__net25 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.28e-6 PS=1.28e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__pm2 n7__i5__i6__i2__net25 n10__i5__clk_buf n8__i5__i6__i2__net22 n328__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i8__pm3 n7__i5__i6__i8__net4 n23__shift n356__vdd n328__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i8__pm5 n12__i5__i6__net35 i5__i6__i8__net4 n9__i5__i6__net34 n328__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i8__pm4 n10__i5__i6__net35 n32__shift n11__i5__r0 n328__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i7__pm3 n7__i5__i6__i7__net4 n10__shift n347__vdd n328__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i7__pm5 n12__i5__i6__net33 i5__i6__i7__net4 n9__i5__i6__net32 n328__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i7__pm4 n10__i5__i6__net33 n19__shift n10__i5__r1 n328__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i6__pm3 n7__i5__i6__i6__net4 n1__shift n338__vdd n328__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i6__pm5 n12__i5__i6__net30 i5__i6__i6__net4 n43__vdd n328__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i6__pm4 n10__i5__i6__net30 n6__shift n3__i5__r2 n328__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__pm1_1__rcx n14__piso_out n5__i4__net1 n368__vdd n328__vdd g45p1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm1 n370__vdd i4__net1 n14__piso_out n328__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi4__pm0 n7__i4__net1 bufin n365__vdd n328__vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi2__pm0_3__rcx n4__piso_outinv n9__piso_out n374__vdd n328__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm0_2__rcx n375__vdd n1__piso_out n4__piso_outinv n328__vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm0_1__rcx n8__piso_outinv n13__piso_out n372__vdd n328__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__pm0 n374__vdd n11__piso_out n8__piso_outinv n328__vdd g45p1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi1__i14__m3_96__rcx n27__vss n22__i1__i14__net1 n133__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_95__rcx n94__chipdriverout n17__i1__i14__net1 n27__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_94__rcx n14__vss n13__i1__i14__net1 n94__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_93__rcx n55__chipdriverout n9__i1__i14__net1 n14__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_92__rcx n1__vss n5__i1__i14__net1 n55__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_91__rcx n16__chipdriverout i1__i14__net1 n1__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=960e-15 AS=960e-15 PD=13.15e-6 PS=13.15e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_90__rcx n66__vss n46__i1__i14__net1 n235__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_89__rcx n196__chipdriverout n41__i1__i14__net1 n66__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_88__rcx n53__vss n38__i1__i14__net1 n196__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_87__rcx n157__chipdriverout n33__i1__i14__net1 n53__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_86__rcx n40__vss n30__i1__i14__net1 n157__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_85__rcx n133__chipdriverout n25__i1__i14__net1 n40__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_84__rcx n105__vss n81__i1__i14__net1 n352__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_83__rcx n313__chipdriverout n77__i1__i14__net1 n105__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_82__rcx n92__vss n66__i1__i14__net1 n313__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_81__rcx n274__chipdriverout n57__i1__i14__net1 n92__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_80__rcx n79__vss n54__i1__i14__net1 n274__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_79__rcx n235__chipdriverout n49__i1__i14__net1 n79__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_78__rcx n144__vss n131__i1__i14__net1 n484__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_77__rcx n430__chipdriverout n125__i1__i14__net1 n144__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_76__rcx n139__vss n113__i1__i14__net1 n430__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_75__rcx n391__chipdriverout n105__i1__i14__net1 n139__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_74__rcx n118__vss n97__i1__i14__net1 n391__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_73__rcx n352__chipdriverout n89__i1__i14__net1 n118__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_72__rcx n183__vss n177__i1__i14__net1 n601__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_71__rcx n580__chipdriverout n173__i1__i14__net1 n183__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_70__rcx n178__vss n161__i1__i14__net1 n580__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_69__rcx n541__chipdriverout n157__i1__i14__net1 n178__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_68__rcx n157__vss n145__i1__i14__net1 n541__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_67__rcx n484__chipdriverout n141__i1__i14__net1 n157__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_66__rcx n230__vss n225__i1__i14__net1 n718__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_65__rcx n679__chipdriverout n217__i1__i14__net1 n230__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_64__rcx n217__vss n209__i1__i14__net1 n679__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_63__rcx n640__chipdriverout n201__i1__i14__net1 n217__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_62__rcx n204__vss n197__i1__i14__net1 n640__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_61__rcx n601__chipdriverout n185__i1__i14__net1 n204__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_60__rcx n261__vss n273__i1__i14__net1 n820__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_59__rcx n781__chipdriverout n269__i1__i14__net1 n261__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_58__rcx n256__vss n257__i1__i14__net1 n781__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_57__rcx n757__chipdriverout n253__i1__i14__net1 n256__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_56__rcx n243__vss n241__i1__i14__net1 n757__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_55__rcx n718__chipdriverout n237__i1__i14__net1 n243__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_54__rcx n308__vss n326__i1__i14__net1 n937__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_53__rcx n898__chipdriverout n313__i1__i14__net1 n308__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_52__rcx n291__vss n306__i1__i14__net1 n898__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_51__rcx n882__chipdriverout n301__i1__i14__net1 n291__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_50__rcx n274__vss n293__i1__i14__net1 n882__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_49__rcx n820__chipdriverout n285__i1__i14__net1 n274__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_48__rcx n937__chipdriverout n333__i1__i14__net1 n321__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_47__rcx n1054__chipdriverout n379__i1__i14__net1 n352__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_46__rcx n347__vss n374__i1__i14__net1 n1054__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_45__rcx n1015__chipdriverout n361__i1__i14__net1 n347__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_44__rcx n334__vss n358__i1__i14__net1 n1015__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_43__rcx n1002__chipdriverout n345__i1__i14__net1 n334__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_42__rcx n321__vss n342__i1__i14__net1 n1002__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_41__rcx n1171__chipdriverout n425__i1__i14__net1 n391__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_40__rcx n386__vss n422__i1__i14__net1 n1171__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_39__rcx n1132__chipdriverout n413__i1__i14__net1 n386__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_38__rcx n373__vss n406__i1__i14__net1 n1132__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_37__rcx n1119__chipdriverout n393__i1__i14__net1 n373__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_36__rcx n352__vss n390__i1__i14__net1 n1119__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_35__rcx n1288__chipdriverout n477__i1__i14__net1 n438__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_34__rcx n417__vss n465__i1__i14__net1 n1288__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_33__rcx n1249__chipdriverout n457__i1__i14__net1 n417__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_32__rcx n404__vss n449__i1__i14__net1 n1249__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_31__rcx n1210__chipdriverout n441__i1__i14__net1 n404__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_30__rcx n391__vss n433__i1__i14__net1 n1210__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_29__rcx n1405__chipdriverout n525__i1__i14__net1 n477__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_28__rcx n456__vss n513__i1__i14__net1 n1405__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_27__rcx n1366__chipdriverout n505__i1__i14__net1 n456__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_26__rcx n443__vss n497__i1__i14__net1 n1366__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_25__rcx n1327__chipdriverout n493__i1__i14__net1 n443__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_24__rcx n438__vss n481__i1__i14__net1 n1327__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_23__rcx n1539__chipdriverout n569__i1__i14__net1 n508__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_22__rcx n503__vss n561__i1__i14__net1 n1539__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_21__rcx n1499__chipdriverout n553__i1__i14__net1 n503__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_20__rcx n482__vss n545__i1__i14__net1 n1499__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_19__rcx n1472__chipdriverout n541__i1__i14__net1 n482__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_18__rcx n477__vss n529__i1__i14__net1 n1472__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_17__rcx n1672__chipdriverout n617__i1__i14__net1 n553__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_16__rcx n534__vss n609__i1__i14__net1 n1672__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_15__rcx n1633__chipdriverout n605__i1__i14__net1 n534__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_14__rcx n521__vss n593__i1__i14__net1 n1633__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_13__rcx n1579__chipdriverout n589__i1__i14__net1 n521__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_12__rcx n508__vss n577__i1__i14__net1 n1579__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_11__rcx n1789__chipdriverout n669__i1__i14__net1 n592__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_10__rcx n587__vss n657__i1__i14__net1 n1789__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_9__rcx n1750__chipdriverout n649__i1__i14__net1 n587__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_8__rcx n566__vss n645__i1__i14__net1 n1750__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_7__rcx n1711__chipdriverout n637__i1__i14__net1 n566__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_6__rcx n553__vss n629__i1__i14__net1 n1711__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_5__rcx n618__vss n705__i1__i14__net1 n1906__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_4__rcx n1867__chipdriverout n701__i1__i14__net1 n618__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_3__rcx n605__vss n689__i1__i14__net1 n1867__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_2__rcx n1823__chipdriverout n685__i1__i14__net1 n605__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3_1__rcx n592__vss n673__i1__i14__net1 n1823__chipdriverout n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m3 n1906__chipdriverout n713__i1__i14__net1 n636__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.15e-6 PS=13.15e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_27__rcx n750__vss n25__i1__net2 n909__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_26__rcx n870__i1__i14__net1 n21__i1__net2 n750__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_25__rcx n729__vss n17__i1__net2 n870__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_24__rcx n831__i1__i14__net1 n13__i1__net2 n729__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_23__rcx n716__vss n10__i1__net2 n831__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_22__rcx n792__i1__i14__net1 n5__i1__net2 n716__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_21__rcx n703__vss n2__i1__net2 n792__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=960e-15 AS=960e-15 PD=13.15e-6 PS=13.15e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_20__rcx n1041__i1__i14__net1 n53__i1__net2 n802__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_19__rcx n781__vss n49__i1__net2 n1041__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_18__rcx n987__i1__i14__net1 n45__i1__net2 n781__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_17__rcx n768__vss n41__i1__net2 n987__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_16__rcx n948__i1__i14__net1 n37__i1__net2 n768__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_15__rcx n755__vss n33__i1__net2 n948__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_14__rcx n909__i1__i14__net1 n29__i1__net2 n755__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_13__rcx n833__vss n105__i1__net2 n1197__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_12__rcx n1143__i1__i14__net1 n101__i1__net2 n833__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_11__rcx n820__vss n93__i1__net2 n1143__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_10__rcx n1104__i1__i14__net1 n85__i1__net2 n820__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_9__rcx n807__vss n73__i1__net2 n1104__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_8__rcx n1098__i1__i14__net1 n65__i1__net2 n807__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_7__rcx n802__vss n57__i1__net2 n1098__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_6__rcx n1325__i1__i14__net1 n181__i1__net2 n908__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.15e-6 PS=13.15e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_5__rcx n880__vss n153__i1__net2 n1325__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_4__rcx n1260__i1__i14__net1 n145__i1__net2 n880__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_3__rcx n859__vss n137__i1__net2 n1260__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_2__rcx n1236__i1__i14__net1 n133__i1__net2 n859__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2_1__rcx n846__vss n121__i1__net2 n1236__i1__i14__net1 n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i14__m2 n1197__i1__i14__net1 n113__i1__net2 n846__vss n1013__vss g45n2svt L=150e-9 W=6.4e-6 AD=1.28e-12 AS=1.28e-12 PD=13.2e-6 PS=13.2e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i11__m0_2__rcx n24__i1__net4 n10__piso_outinv n1621__vss n1013__vss g45n2svt L=150e-9 W=640e-9 AD=96e-15 AS=96e-15 PD=1.63e-6 PS=1.63e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i11__m1_2__rcx n5__i1__i11__outinv n27__piso_out n1622__vss n1013__vss g45n2svt L=150e-9 W=640e-9 AD=128e-15 AS=128e-15 PD=1.63e-6 PS=1.63e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i11__m1_1__rcx n1623__vss n25__piso_out n5__i1__i11__outinv n1013__vss g45n2svt L=150e-9 W=640e-9 AD=128e-15 AS=128e-15 PD=1.68e-6 PS=1.68e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i11__m1 n9__i1__i11__outinv n22__piso_out n1623__vss n1013__vss g45n2svt L=150e-9 W=640e-9 AD=96e-15 AS=96e-15 PD=1.63e-6 PS=1.63e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i11__m0_1__rcx n1621__vss n12__piso_outinv n27__i1__net4 n1013__vss g45n2svt L=150e-9 W=640e-9 AD=128e-15 AS=128e-15 PD=1.68e-6 PS=1.68e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i11__m0 n27__i1__net4 n14__piso_outinv n1613__vss n1013__vss g45n2svt L=150e-9 W=640e-9 AD=128e-15 AS=128e-15 PD=1.63e-6 PS=1.63e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_20__rcx n262__i1__net2 n28__i1__i13__net1 n1553__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_19__rcx n1307__vss n23__i1__i13__net1 n262__i1__net2 n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_18__rcx n253__i1__net2 n19__i1__i13__net1 n1307__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_17__rcx n1300__vss n15__i1__i13__net1 n253__i1__net2 n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_16__rcx n239__i1__net2 n11__i1__i13__net1 n1300__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_15__rcx n1293__vss n7__i1__i13__net1 n239__i1__net2 n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_14__rcx n235__i1__net2 n3__i1__i13__net1 n1293__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=384e-15 AS=384e-15 PD=5.47e-6 PS=5.47e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_13__rcx n1553__vss n31__i1__i13__net1 n271__i1__net2 n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_12__rcx n298__i1__net2 n60__i1__i13__net1 n1594__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_11__rcx n1588__vss n55__i1__i13__net1 n298__i1__net2 n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_10__rcx n289__i1__net2 n52__i1__i13__net1 n1588__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_9__rcx n1567__vss n47__i1__i13__net1 n289__i1__net2 n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_8__rcx n280__i1__net2 n44__i1__i13__net1 n1567__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_7__rcx n1561__vss n39__i1__i13__net1 n280__i1__net2 n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_6__rcx n271__i1__net2 n36__i1__i13__net1 n1561__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_5__rcx n320__i1__net2 n124__i1__i13__net1 n1625__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.47e-6 PS=5.47e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_4__rcx n1608__vss n99__i1__i13__net1 n320__i1__net2 n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_3__rcx n311__i1__net2 n92__i1__i13__net1 n1608__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_2__rcx n1602__vss n83__i1__i13__net1 n311__i1__net2 n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1_1__rcx n307__i1__net2 n80__i1__i13__net1 n1602__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m1 n1594__vss n67__i1__i13__net1 n307__i1__net2 n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m0_5__rcx n181__i1__i13__net1 n50__i1__net3 n1650__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.47e-6 PS=5.47e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m0_4__rcx n1645__vss n46__i1__net3 n181__i1__i13__net1 n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m0_3__rcx n170__i1__i13__net1 n42__i1__net3 n1645__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m0_2__rcx n1639__vss n38__i1__net3 n170__i1__i13__net1 n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m0_1__rcx n159__i1__i13__net1 n34__i1__net3 n1639__vss n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=512e-15 AS=512e-15 PD=5.52e-6 PS=5.52e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i13__m0 n1631__vss n30__i1__net3 n159__i1__i13__net1 n1013__vss g45n2svt L=150e-9 W=2.56e-6 AD=384e-15 AS=384e-15 PD=5.47e-6 PS=5.47e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m2_1__rcx n66__i1__i12__net1 n5__i1__net4 n1572__vss n1013__vss g45n2svt L=150e-9 W=640e-9 AD=128e-15 AS=128e-15 PD=1.63e-6 PS=1.63e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m2 n1580__vss i1__net4 n66__i1__i12__net1 n1013__vss g45n2svt L=150e-9 W=640e-9 AD=96e-15 AS=96e-15 PD=1.63e-6 PS=1.63e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m3_6__rcx n29__i1__net3 n25__i1__i12__net1 n1581__vss n1013__vss g45n2svt L=150e-9 W=640e-9 AD=128e-15 AS=128e-15 PD=1.63e-6 PS=1.63e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m3_5__rcx n1582__vss n21__i1__i12__net1 n29__i1__net3 n1013__vss g45n2svt L=150e-9 W=640e-9 AD=128e-15 AS=128e-15 PD=1.68e-6 PS=1.68e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m3_4__rcx n16__i1__net3 n17__i1__i12__net1 n1582__vss n1013__vss g45n2svt L=150e-9 W=640e-9 AD=128e-15 AS=128e-15 PD=1.68e-6 PS=1.68e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m3_3__rcx n1583__vss n13__i1__i12__net1 n16__i1__net3 n1013__vss g45n2svt L=150e-9 W=640e-9 AD=128e-15 AS=128e-15 PD=1.68e-6 PS=1.68e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m3_2__rcx n9__i1__net3 n9__i1__i12__net1 n1583__vss n1013__vss g45n2svt L=150e-9 W=640e-9 AD=128e-15 AS=128e-15 PD=1.68e-6 PS=1.68e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m3_1__rcx n1579__vss n5__i1__i12__net1 n9__i1__net3 n1013__vss g45n2svt L=150e-9 W=640e-9 AD=128e-15 AS=128e-15 PD=1.68e-6 PS=1.68e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi1__i12__m3 n2__i1__net3 i1__i12__net1 n1579__vss n1013__vss g45n2svt L=150e-9 W=640e-9 AD=96e-15 AS=96e-15 PD=1.63e-6 PS=1.63e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
mi5__i8__i5__nm0_2__rcx n17__i5__i8__net5 n84__i5__clk4 n1198__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i5__nm0_1__rcx n16__i5__i8__net5 n81__i5__clk4 n1199__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i5__nm0 n1198__vss n83__i5__clk4 n16__i5__i8__net5 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i4__nm0_2__rcx n22__i5__i8__net1 n9__i5__i8__net2 n1210__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i4__nm0_1__rcx n21__i5__i8__net1 n6__i5__i8__net2 n1211__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i4__nm0 n1210__vss n8__i5__i8__net2 n21__i5__i8__net1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i6__nm0_2__rcx n13__i5__i8__net4 n26__i5__clk_buf n1221__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i6__nm0_1__rcx n11__i5__i8__net4 n23__i5__clk_buf n1222__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i6__nm0 n1221__vss n25__i5__clk_buf n11__i5__i8__net4 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__nm3_1__rcx n1208__vss n5__i5__i8__i10__net22 i5__i8__i10__net23 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__nm3 n4__i5__i8__i10__net23 n7__i5__i8__i10__net22 n1208__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__nm2_1__rcx n93__i5__clk4 n14__i5__i8__net2 n4__i5__i8__i10__net23 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__nm2 n7__i5__i8__i10__net23 n13__i5__i8__net2 n93__i5__clk4 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__nm4_1__rcx n1207__vss n63__reset n96__i5__clk4 n1013__vss g45n1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__nm4 n95__i5__clk4 n60__reset n1207__vss n1013__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__nm1_1__rcx n1209__vss n5__i5__i8__net5 i5__i8__i10__net21 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__nm1 n4__i5__i8__i10__net21 n7__i5__i8__net5 n1209__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__nm0_1__rcx n10__i5__i8__i10__net22 n14__i5__i8__net1 n4__i5__i8__i10__net21 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i10__nm0 n8__i5__i8__i10__net21 n11__i5__i8__net1 n10__i5__i8__i10__net22 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__nm3_1__rcx n1219__vss n5__i5__i8__i9__net22 i5__i8__i9__net23 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__nm3 n4__i5__i8__i9__net23 n7__i5__i8__i9__net22 n1219__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__nm2_1__rcx n25__i5__i8__net2 n41__i5__clk_buf n4__i5__i8__i9__net23 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__nm2 n8__i5__i8__i9__net23 n40__i5__clk_buf n25__i5__i8__net2 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__nm4_1__rcx n1218__vss n50__reset n28__i5__i8__net2 n1013__vss g45n1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__nm4 n26__i5__i8__net2 n47__reset n1218__vss n1013__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__nm1_1__rcx n1220__vss n5__i5__i8__net1 i5__i8__i9__net21 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__nm1 n4__i5__i8__i9__net21 n7__i5__i8__net1 n1220__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__nm0_1__rcx n10__i5__i8__i9__net22 n4__i5__i8__net4 n4__i5__i8__i9__net21 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i9__nm0 n7__i5__i8__i9__net21 i5__i8__net4 n10__i5__i8__i9__net22 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i8__nm2 n46__shift n3__i5__i8__i8__net1 n1195__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i8__nm1 n6__i5__i8__i8__net1 n88__i5__clk4 n1197__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i8__i8__nm0 n1196__vss n31__i5__i8__net2 n6__i5__i8__i8__net1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i2__nm3 n2__i5__i7__i1__i2__net25 n4__i5__i7__i1__i2__net22 n1281__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i2__nm2 n10__i5__i7__y3out n56__i5__clk4 i5__i7__i1__i2__net25 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i2__nm4 n6__i5__i7__y3out n26__reset n1280__vss n1013__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i2__nm1 n2__i5__i7__i1__i2__net23 n4__y3 n1282__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i2__nm0 n7__i5__i7__i1__i2__net22 n21__i5__i7__i1__net1 i5__i7__i1__i2__net23 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i1__nm3 n2__i5__i7__i1__i1__net25 n4__i5__i7__i1__i1__net22 n1284__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i1__nm2 n8__i5__i7__y2out n42__i5__clk4 i5__i7__i1__i1__net25 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i1__nm4 n4__i5__i7__y2out n18__reset n1283__vss n1013__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i1__nm1 n2__i5__i7__i1__i1__net23 n4__y2 n1285__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i1__nm0 n7__i5__i7__i1__i1__net22 n16__i5__i7__i1__net1 i5__i7__i1__i1__net23 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i0__nm3 n2__i5__i7__i1__i0__net25 n4__i5__i7__i1__i0__net22 n1287__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i0__nm2 n5__i5__i7__y1out n28__i5__clk4 i5__i7__i1__i0__net25 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i0__nm4 i5__i7__y1out n7__reset n1286__vss n1013__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i0__nm1 n2__i5__i7__i1__i0__net23 n4__y1 n1288__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i0__nm0 n7__i5__i7__i1__i0__net22 n5__i5__i7__i1__net1 i5__i7__i1__i0__net23 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i3__nm3 n2__i5__i7__i1__i3__net25 n4__i5__i7__i1__i3__net22 n1290__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i3__nm2 n5__i5__i7__y0out n13__i5__clk4 i5__i7__i1__i3__net25 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i3__nm4 i5__i7__y0out n3__reset n1289__vss n1013__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i3__nm1 n2__i5__i7__i1__i3__net23 n4__y0 n1291__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i3__nm0 n7__i5__i7__i1__i3__net22 i5__i7__i1__net1 i5__i7__i1__i3__net23 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i1__i4__nm0 n8__i5__i7__i1__net1 n6__i5__clk4 n1267__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i2__nm3 n2__i5__i7__i0__i2__net25 n4__i5__i7__i0__i2__net22 n1092__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i2__nm2 n8__i5__i7__x3out n54__i5__clk4 i5__i7__i0__i2__net25 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i2__nm4 n4__i5__i7__x3out n24__reset n1094__vss n1013__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i2__nm1 n2__i5__i7__i0__i2__net23 n4__x3 n1090__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i2__nm0 n7__i5__i7__i0__i2__net22 n21__i5__i7__i0__net1 i5__i7__i0__i2__net23 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i1__nm3 n2__i5__i7__i0__i1__net25 n4__i5__i7__i0__i1__net22 n1083__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i1__nm2 n8__i5__i7__x2out n40__i5__clk4 i5__i7__i0__i1__net25 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i1__nm4 n4__i5__i7__x2out n16__reset n1085__vss n1013__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i1__nm1 n2__i5__i7__i0__i1__net23 n4__x2 n1081__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i1__nm0 n7__i5__i7__i0__i1__net22 n16__i5__i7__i0__net1 i5__i7__i0__i1__net23 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i0__nm3 n2__i5__i7__i0__i0__net25 n4__i5__i7__i0__i0__net22 n1074__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i0__nm2 n5__i5__i7__x1out n26__i5__clk4 i5__i7__i0__i0__net25 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i0__nm4 i5__i7__x1out n5__reset n1076__vss n1013__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i0__nm1 n2__i5__i7__i0__i0__net23 n4__x1 n1069__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i0__nm0 n7__i5__i7__i0__i0__net22 n5__i5__i7__i0__net1 i5__i7__i0__i0__net23 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i3__nm3 n2__i5__i7__i0__i3__net25 n4__i5__i7__i0__i3__net22 n1071__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i3__nm2 n5__i5__i7__x0out n11__i5__clk4 i5__i7__i0__i3__net25 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i3__nm4 i5__i7__x0out n1__reset n1070__vss n1013__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i3__nm1 n2__i5__i7__i0__i3__net23 n4__x0 n1072__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i3__nm0 n7__i5__i7__i0__i3__net22 i5__i7__i0__net1 i5__i7__i0__i3__net23 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i0__i4__nm0 n8__i5__i7__i0__net1 n3__i5__clk4 n1067__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i5__i0__nm0 n12__i5__i7__xor3 n12__i5__i7__xor2 n9__i5__i7__net47 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=23.4e-15 AS=23.4e-15 PD=830e-9 PS=830e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i5__i0__nm1 n9__i5__i7__net47 n4__i5__i7__i5__net1 n1276__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=47.4e-15 AS=47.4e-15 PD=835e-9 PS=835e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i5__i1__nm0 n26__i5__i7__xor3 n5__i5__i7__i5__net1 n11__i5__i7__net51 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=27e-15 AS=27e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i5__i1__nm1 n11__i5__i7__net51 n3__i5__i7__xor3 n13__i5__i7__i5__net1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=66.6e-15 AS=66.6e-15 PD=1.025e-6 PS=1.025e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i5__i2__nm0 n9__i5__i7__i5__net1 n3__i5__i7__xor2 n1277__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i6__i0__nm0 n12__i5__i7__net50 n5__i5__i7__net51 n7__i5__i7__net46 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=23.4e-15 AS=23.4e-15 PD=830e-9 PS=830e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i6__i0__nm1 n7__i5__i7__net46 n4__i5__i7__i6__net1 n1123__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=47.4e-15 AS=47.4e-15 PD=835e-9 PS=835e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i6__i1__nm0 n24__i5__i7__net50 n5__i5__i7__i6__net1 n7__i5__r0 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=27e-15 AS=27e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i6__i1__nm1 n7__i5__r0 n3__i5__i7__net50 n13__i5__i7__i6__net1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=66.6e-15 AS=66.6e-15 PD=1.025e-6 PS=1.025e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i6__i2__nm0 n11__i5__i7__i6__net1 n3__i5__i7__net51 n1120__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i4__i0__nm0 n12__i5__i7__xor0 n12__i5__i7__xor1 n7__i5__i7__net44 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=23.4e-15 AS=23.4e-15 PD=830e-9 PS=830e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i4__i0__nm1 n7__i5__i7__net44 n4__i5__i7__i4__net1 n1114__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=47.4e-15 AS=47.4e-15 PD=835e-9 PS=835e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i4__i1__nm0 n26__i5__i7__xor0 n5__i5__i7__i4__net1 n7__i5__i7__net50 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=27e-15 AS=27e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i4__i1__nm1 n7__i5__i7__net50 n3__i5__i7__xor0 n13__i5__i7__i4__net1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=66.6e-15 AS=66.6e-15 PD=1.025e-6 PS=1.025e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i4__i2__nm0 n9__i5__i7__i4__net1 n3__i5__i7__xor1 n1111__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i1__i0__nm0 n17__i5__i7__net46 i5__i7__i7__i1__net1 n4__i5__r1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=27e-15 AS=27e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i1__i0__nm1 n4__i5__r1 n3__i5__i7__net46 n6__i5__i7__i7__i1__net1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=66.6e-15 AS=66.6e-15 PD=1.025e-6 PS=1.025e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i1__i1__nm0 n4__i5__i7__i7__i1__net1 n3__i5__i7__i7__net1 n1274__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i0__i0__nm0 n17__i5__i7__net44 i5__i7__i7__i0__net1 n12__i5__i7__i7__net1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=27e-15 AS=27e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i0__i0__nm1 n12__i5__i7__i7__net1 n3__i5__i7__net44 n6__i5__i7__i7__i0__net1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=66.6e-15 AS=66.6e-15 PD=1.025e-6 PS=1.025e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i0__i1__nm0 n4__i5__i7__i7__i0__net1 n3__i5__i7__net47 n1275__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i4__nm3 i5__i7__i7__i4__net4 n10__i5__i7__net44 n1272__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=37.8e-15 AS=37.8e-15 PD=765e-9 PS=765e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i4__nm2 n5__i5__i7__i7__net3 n3__i5__i7__i7__net2 i5__i7__i7__i4__net4 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=37.8e-15 AS=37.8e-15 PD=870e-9 PS=870e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i4__nm0 i5__i7__i7__i4__net1 n11__i5__i7__net46 n5__i5__i7__i7__net3 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=37.8e-15 AS=37.8e-15 PD=870e-9 PS=870e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i4__nm1 n1271__vss n18__i5__i7__i7__net1 i5__i7__i7__i4__net1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=27e-15 AS=27e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i2__nm0 n7__i5__i7__i7__net2 n8__i5__i7__i7__net1 n1273__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i7__i3__nm0 n11__i5__r2 n3__i5__i7__i7__net3 n1270__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i9__i0__nm0 n17__i5__i7__x3out i5__i7__i9__net1 n7__i5__i7__xor3 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=27e-15 AS=27e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i9__i0__nm1 n7__i5__i7__xor3 n3__i5__i7__x3out n6__i5__i7__i9__net1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=66.6e-15 AS=66.6e-15 PD=1.025e-6 PS=1.025e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i9__i1__nm0 n4__i5__i7__i9__net1 n3__i5__i7__y3out n1278__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i8__i0__nm0 n17__i5__i7__x2out i5__i7__i8__net1 n7__i5__i7__xor2 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=27e-15 AS=27e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i8__i0__nm1 n7__i5__i7__xor2 n3__i5__i7__x2out n6__i5__i7__i8__net1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=66.6e-15 AS=66.6e-15 PD=1.025e-6 PS=1.025e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i8__i1__nm0 n4__i5__i7__i8__net1 n3__i5__i7__y2out n1279__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i2__i0__nm0 n17__i5__i7__x0out i5__i7__i2__net1 n7__i5__i7__xor0 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=27e-15 AS=27e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i2__i0__nm1 n7__i5__i7__xor0 n10__i5__i7__x0out n6__i5__i7__i2__net1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=66.6e-15 AS=66.6e-15 PD=1.025e-6 PS=1.025e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i2__i1__nm0 n4__i5__i7__i2__net1 n10__i5__i7__y0out n1105__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i3__i0__nm0 n17__i5__i7__x1out i5__i7__i3__net1 n7__i5__i7__xor1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=27e-15 AS=27e-15 PD=1.02e-6 PS=1.02e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i3__i0__nm1 n7__i5__i7__xor1 n10__i5__i7__x1out n6__i5__i7__i3__net1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=66.6e-15 AS=66.6e-15 PD=1.025e-6 PS=1.025e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i7__i3__i1__nm0 n4__i5__i7__i3__net1 n10__i5__i7__y1out n1099__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i9__nm1_3__rcx n699__vss n17__i5__i9__net21 n48__i5__clk_buf n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i9__nm0_1__rcx n20__i5__i9__net21 n3__clk_out n1269__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i9__nm0 n1268__vss n2__clk_out n20__i5__i9__net21 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i9__nm1_2__rcx n47__i5__clk_buf n4__i5__i9__net21 n631__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i9__nm1_1__rcx n635__vss n9__i5__i9__net21 n47__i5__clk_buf n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i9__nm1 n48__i5__clk_buf n13__i5__i9__net21 n635__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i9__nm0_2__rcx n13__i5__i6__net31 n9__i5__clk_buf n1132__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i9__nm0_1__rcx n11__i5__i6__net31 n6__i5__clk_buf n1129__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i9__nm0 n1132__vss n8__i5__clk_buf n11__i5__i6__net31 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__nm3_1__rcx n1170__vss n5__i5__i6__i5__net22 i5__i6__i5__net23 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__nm3 n4__i5__i6__i5__net23 n7__i5__i6__i5__net22 n1170__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__nm2_1__rcx n8__bufin n61__i5__clk_buf n4__i5__i6__i5__net23 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__nm2 n8__i5__i6__i5__net23 n60__i5__clk_buf n8__bufin n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__nm4_1__rcx n1172__vss n59__reset n9__bufin n1013__vss g45n1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__nm4 n4__bufin n56__reset n1172__vss n1013__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__nm1_1__rcx n1165__vss n5__i5__i6__net35 i5__i6__i5__net21 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__nm1 n4__i5__i6__i5__net21 n7__i5__i6__net35 n1165__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__nm0_1__rcx n10__i5__i6__i5__net22 n35__i5__i6__net31 n4__i5__i6__i5__net21 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i5__nm0 n8__i5__i6__i5__net21 n32__i5__i6__net31 n10__i5__i6__i5__net22 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__nm3_1__rcx n1156__vss n5__i5__i6__i4__net22 i5__i6__i4__net23 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__nm3 n4__i5__i6__i4__net23 n7__i5__i6__i4__net22 n1156__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__nm2_1__rcx n5__i5__i6__net34 n38__i5__clk_buf n4__i5__i6__i4__net23 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__nm2 n7__i5__i6__i4__net23 n37__i5__clk_buf n5__i5__i6__net34 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__nm4_1__rcx n1158__vss n46__reset n6__i5__i6__net34 n1013__vss g45n1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__nm4 i5__i6__net34 n43__reset n1158__vss n1013__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__nm1_1__rcx n1153__vss n5__i5__i6__net33 i5__i6__i4__net21 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__nm1 n4__i5__i6__i4__net21 n7__i5__i6__net33 n1153__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__nm0_1__rcx n10__i5__i6__i4__net22 n21__i5__i6__net31 n4__i5__i6__i4__net21 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i4__nm0 n7__i5__i6__i4__net21 n18__i5__i6__net31 n10__i5__i6__i4__net22 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__nm3_1__rcx n1142__vss n5__i5__i6__i2__net22 i5__i6__i2__net23 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__nm3 n4__i5__i6__i2__net23 n7__i5__i6__i2__net22 n1142__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__nm2_1__rcx n5__i5__i6__net32 n14__i5__clk_buf n4__i5__i6__i2__net23 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__nm2 n7__i5__i6__i2__net23 n13__i5__clk_buf n5__i5__i6__net32 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__nm4_1__rcx n1144__vss n39__reset n6__i5__i6__net32 n1013__vss g45n1svt L=45e-9 W=480e-9 AD=76.8e-15 AS=76.8e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__nm4 i5__i6__net32 n36__reset n1144__vss n1013__vss g45n1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.26e-6 PS=1.26e-6 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__nm1_1__rcx n1139__vss n5__i5__i6__net30 i5__i6__i2__net21 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__nm1 n4__i5__i6__i2__net21 n7__i5__i6__net30 n1139__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__nm0_1__rcx n10__i5__i6__i2__net22 n4__i5__i6__net31 n4__i5__i6__i2__net21 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=800e-9 PS=800e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i2__nm0 n7__i5__i6__i2__net21 i5__i6__net31 n10__i5__i6__i2__net22 n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i8__nm3 n5__i5__i6__i8__net4 n25__shift n1162__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i8__nm5 n14__i5__i6__net35 n30__shift n10__i5__i6__net34 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i8__nm6 n8__i5__i6__net35 n3__i5__i6__i8__net4 n13__i5__r0 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i7__nm3 n5__i5__i6__i7__net4 n12__shift n1146__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i7__nm5 n14__i5__i6__net33 n17__shift n10__i5__i6__net32 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i7__nm6 n8__i5__i6__net33 n3__i5__i6__i7__net4 n12__i5__r1 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i6__nm3 n5__i5__i6__i6__net4 n3__shift n1134__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i6__nm5 n14__i5__i6__net30 n4__shift n45__vdd n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi5__i6__i6__nm6 n8__i5__i6__net30 n3__i5__i6__i6__net4 n5__i5__r2 n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm1_1__rcx n17__piso_out n3__i4__net1 n1179__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=38.4e-15 AS=38.4e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm1 n1181__vss n2__i4__net1 n17__piso_out n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=780e-9 PS=780e-9 NRD=1.16667 NRS=1.16667 M=1
mi4__nm0 n9__i4__net1 n3__bufin n1176__vss n1013__vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm0_3__rcx n7__piso_outinv n8__piso_out n1193__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm0_2__rcx n1194__vss n7__piso_out n7__piso_outinv n1013__vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm0_1__rcx n6__piso_outinv n12__piso_out n1184__vss n1013__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=540e-9 PS=540e-9 NRD=1.16667 NRS=1.16667 M=1
mi2__nm0 n1193__vss n10__piso_out n6__piso_outinv n1013__vss g45n1svt L=45e-9 W=120e-9 AD=19.2e-15 AS=19.2e-15 PD=560e-9 PS=560e-9 NRD=1.16667 NRS=1.16667 M=1
.END
