** Generated for: hspiceD
** Generated on: Dec 2, 2024
** Design library name: final_project
** Design cell name: Adder_Comp
** Design view name: schematic

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Subcircuit Definitions

** Pass-Transistor Logic XOR Gate
.subckt ptl_Xor a b bnot out vdd vss
mnm1 out a bnot vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0 a bnot out vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm1 out a b vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm0 a b out vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
.ends ptl_Xor

** Inverter
.subckt inv_n120 d q vdd vss
mpm0 q d vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm0 q d vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
.ends inv_n120

** XOR Gate
.subckt XOR a b out vdd vss
xi0 a b net1 out vdd vss ptl_Xor
xi1 b net1 vdd vss inv_n120
.ends XOR

** AND
** AND Gate
.subckt AND a b bnot out vdd vss
mnm1 out bnot vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0 a b out vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm0 out bnot a vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
.ends AND

** Half Adder
.subckt HalfAdder a b cout s vdd vss
xi0 a b net1 cout vdd vss AND
xi1 a b net1 s vdd vss ptl_Xor
xi2 b net1 vdd vss inv_n120
.ends HalfAdder

** Cout Logic
.subckt CoutLogic a coutnot cin p pnot vdd vss
mpm3 coutnot p net3 vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm2 net3 a vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm1 coutnot cin net2 vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm0 net2 pnot vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm3 net4 a vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm2 coutnot pnot net4 vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm1 net1 p vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0 coutnot cin net1 vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
.ends CoutLogic

** Full Adder
.subckt FullAdder a b cin cout s vdd vss
xi1 cin net1 s vdd vss XOR
xi0 a b net1 vdd vss XOR
xi3 net3 cout vdd vss inv_n120
xi2 net1 net2 vdd vss inv_n120
xi4 a net3 cin net1 net2 vdd vss CoutLogic
.ends FullAdder

** Adder_Comp
.subckt Adder_Comp x0 x1 x2 x3 y0 y1 y2 y3 r0 r1 r2 vdd vss
xi3 x3 y3 net3 vdd vss XOR
xi2 x2 y2 net4 vdd vss XOR
xi1 x1 y1 net2 vdd vss XOR
xi0 x0 y0 net1 vdd vss XOR
xi6 net5 net6 net9 r0 vdd vss HalfAdder
xi5 net3 net4 net8 net6 vdd vss HalfAdder
xi4 net1 net2 net10 net5 vdd vss HalfAdder
xi7 net8 net10 net9 r2 r1 vdd vss FullAdder
.ends Adder_Comp

** Testbench
.lib '/class/ece482/gpdk045_mos' TT

** Simulation parameters
.param TCK = 0.4167n
.param trf_ck = 5p
.param CK_pw = 0.5*TCK
.param sim_end = 50*TCK
.param trf_ip_reset = 50p
.param reset_delay = 0
.param reset_delay2 = 25*TCK
.param reset_pw = 0.9n
.param reset_pw2 = 3n
.param input_delay = 0.5n
.param input_pw = 4*TCK

** Clock signals
vCK CK 0 pulse(0 1.1 0 5p 5p 0.5*TCK TCK)

** Input signals
** X Inputs: Binary sequences with specific delays
vX3 x3 0 PWL(
+   0 0
+   input_delay 0
+   input_delay+input_pw 1.1
+   input_delay+2*input_pw 0
+   input_delay+3*input_pw 1.1
+   sim_end 0)

vX2 x2 0 PWL(
+   0 0
+   input_delay 0
+   input_delay+input_pw 1.1
+   input_delay+2*input_pw 1.1
+   input_delay+3*input_pw 0
+   sim_end 0)

vX1 x1 0 PWL(
+   0 0
+   input_delay 0
+   input_delay+input_pw 0
+   input_delay+2*input_pw 1.1
+   input_delay+3*input_pw 0
+   sim_end 0)

vX0 x0 0 PWL(
+   0 0
+   input_delay 0
+   input_delay+input_pw 1.1
+   input_delay+2*input_pw 0
+   input_delay+3*input_pw 0
+   sim_end 1.1)

** Y Inputs: Binary sequences with specific delays
vY3 y3 0 PWL(
+   0 0
+   input_delay 0
+   input_delay+input_pw 0
+   input_delay+2*input_pw 0
+   input_delay+3*input_pw 1.1
+   sim_end 1.1)

vY2 y2 0 PWL(
+   0 0
+   input_delay 0
+   input_delay+input_pw 1.1
+   sim_end 1.1)

vY1 y1 0 PWL(
+   0 0
+   input_delay 0
+   input_delay+input_pw 1.1
+   input_delay+2*input_pw 1.1
+   input_delay+3*input_pw 0
+   sim_end 0)

vY0 y0 0 PWL(
+   0 0
+   sim_end 0)


** Power supplies
vVDD VDD 0 1.1
vVSS VSS 0 0

** Circuit instantiation
xi0 x0 x1 x2 x3 y0 y1 y2 y3 r0 r1 r2 VDD VSS Adder_Comp

** Transient analysis
.tran 0 sim_end

.option post
.end
